// file name: parameters.vh	
//constants
`define w	64
`define b	8
`define L	0
`define r	168 // max default value of r (40+512/4)
`define n 	89
`define c 	16

//IV 

`define V0          64'h0000000000000000
`define V1          64'h0000000000000000
`define V2          64'h0000000000000000
`define V3          64'h0000000000000000
`define V4          64'h0000000000000000
`define V5          64'h0000000000000000
`define V6          64'h0000000000000000
`define V7          64'h0000000000000000
`define V8          64'h0000000000000000
`define V9          64'h0000000000000000
`define V10         64'h0000000000000000
`define V11         64'h0000000000000000
`define V12         64'h0000000000000000
`define V13         64'h0000000000000000
`define V14         64'h0000000000000000
`define V15         64'h0000000000000000

`define IV			{`V15	,`V14	,`V13	,`V12	,`V11	,`V10	,`V9	,`V8	,`V7	,`V6	,`V5	,`V4	,`V3	,`V2	,`V1	,`V0}

//Q vector
`define	Q0 			64'h7311c2812425cfa0
`define	Q1 			64'h6432286434aac8e7
`define	Q2 			64'hb60450e9ef68b7c1
`define	Q3 			64'he8fb23908d9f06f1
`define	Q4 			64'hdd2e76cba691e5bf
`define	Q5 			64'h0cd0d63b2c30bc41
`define	Q6 			64'h1f8ccf6823058f8a
`define	Q7 			64'h54e5ed5b88e3775d
`define	Q8 			64'h4ad12aae0a6d6031
`define	Q9 			64'h3e7f16bb88222e0d
`define	Q10 		64'h8af8671d3fb50c2c
`define	Q11			64'h995ad1178bd25c31
`define	Q12			64'hc878c1dd04c4b633
`define	Q13 		64'h3b72066c7a1552ac
`define	Q14 		64'h0d6f3522631effcb
 
 //Q_array[15*w-1:0]
`define Q_array     {`Q14,`Q13,`Q12,`Q11,`Q10,`Q9,`Q8,`Q7,`Q6,`Q5,`Q4,`Q3,`Q2,`Q1,`Q0}

//S vector
/*  S_0^'=64'h123456789abcdef
	S^*=64'h7311c2812425cfa0
	S_(j+1)^'=(S_j^'<< 1)?(S_j^' and S^* ) */

`define	S0 			64'h0123456789abcdef
`define	S1 			64'h0347cace1376567e
`define	S2 			64'h058e571c26c8eadc
`define	S3 			64'h0a1cec3869911f38
`define	S4 			64'h16291870f3233150
`define	S5 			64'h3e5330e1c66763a0
`define	S6 			64'h4eb7614288eb84e0
`define	S7 			64'hdf7f828511f68d60
`define	S8 			64'hedee878b23c997e1
`define	S9 			64'hbadd8d976792a863
`define	S10 		64'h47aa9bafeb25d8e7
`define	S11			64'hcc55b5def66e796e
`define	S12			64'hd8baeb3dc8f8bbfd
`define	S13 		64'he165147a91d1fc5b
`define	S14 		64'ha3cb28f523a234b7
`define	S15 		64'h6497516b67646dcf
`define	S16 		64'ha93fe2d7eaec961e
`define	S17			64'h736e072ef5fdaa3d
`define	S18 		64'h95dc0c5dcfdede5a
`define	S19			64'h3aa818ba9bb972b5
`define	S20			64'h475031f53753a7ca
`define	S21 		64'hcdb0636b4aa6c814
`define	S22 		64'hda7084d795695829
`define	S23			64'he6f1892e2ef3f873
`define	S24			64'haff2925c79c638c7
`define	S25 		64'h7cf5a6b8d388790f
`define	S26			64'h89facff1a710bb1e
`define	S27			64'h12e55d626a21fd3d
`define	S28 		64'h37cbfac4f462375a
`define	S29 		64'h5c963709cce469b4	
`define S30 		64'he93c6c129dec9ac8
`define S31 		64'hb36898253ffdbf11
`define	S32 		64'h55d1b04b5bdef123
`define	S33 		64'hfab2e097b7b92366
`define	S34 		64'h877501ae4b5345ed
`define	S35 		64'h0dfb03dc96a7ce7b
`define	S36 		64'h1ae70539296a52d6
`define	S37 		64'h27cf0a7372f4e72c
`define	S38 		64'h6c9f16e7c5cd0978
`define	S39 		64'hb92f2f4e8f9f1bd0
`define	S40 		64'h435f5c9d1b3b3c21
`define	S41 		64'hc5aff9bb36577462
`define	S42 		64'hca5e33f748abace5
`define	S43 		64'hd6ac656f9176d56b
`define	S44 		64'hff588ade22c96ff7
`define	S45 		64'h8da1973c6593904f
`define	S46 		64'h1a42ac78ef26a09f
`define	S47 		64'h2685d8f1fa69c1be
`define	S48 		64'h6f0a7162d4f242dc
`define	S49 		64'hbd14a2c5adc4c738
`define	S50 		64'h4b39c70a7f8d4951
`define	S51 		64'hd5624c14db1fdba2
`define	S52 		64'hfbc4d829b63a7ce5
`define	S53 		64'h848970524854b56b
`define	S54 		64'h0913a0a490adeff7
`define	S55 		64'h1336c1c9217e104e
`define	S56 		64'h357d431362d8209c
`define	S57 		64'h5bebc427e5b041b8
`define	S58 		64'he4d6484eef40c2d0
`define	S59 		64'ha9bcd09dfa814721
`define	S60 		64'h726961bad503c963
`define	S61 		64'h96d383f5ae065be6
`define	S62 		64'h3fb6856a7808fc6d
`define	S63 		64'h4c7d8ad4d01134fa
`define	S64 		64'hd8ea9729a0236d54
`define	S65 		64'he1d5ac52606797a9
`define	S66 		64'ha2bad8a4e0eaa8f3
`define	S67 		64'h676571c9e1f5d947
`define	S68 		64'hadcba312e3ce7b8e
`define	S69 		64'h7a96c425e798bc9d
`define	S70 		64'h873d484aeb31f5ba
`define	S71 		64'h0d6bd095f6422ed5
`define	S72 		64'h1bd661aac884532a
`define	S73 		64'h24bc83d5910ce574
`define	S74 		64'h6969852a221d0fc8
`define	S75 		64'hb3d28a54643f1010
`define	S76 		64'h54b596a8ec5b2021
`define	S77 		64'hf97aafd1fcb74062
`define	S78 		64'h83e5dd22dd4bc0e5
`define	S79 		64'h04ca7a45be96416b
`define	S80 		64'h0994b68a5928c3f6
`define	S81 		64'h1239ef94b271444c
`define	S82 		64'h36621da944c3cc98
`define	S83 		64'h5ec43bd38d8655b0
`define	S84 		64'hef8875261f08eec0
`define	S85 		64'hbc10aa4c3a111301
`define	S86 		64'h4831d69854232503
`define	S87 		64'hd0726fb0ac674f06
`define	S88 		64'hf0f49de17cebd10d
`define	S89 		64'h91f9bb43ddf6631b
`define	S90 		64'h32e2f486bfc88537
`define	S91 		64'h57c5298d5b918f4e
`define	S92 		64'hfc8b539bb722919c
`define	S93 		64'h8917e5b64a65a2b9
`define	S94 		64'h133e0bec94eec7d3
`define	S95 		64'h356c15592df94826
`define	S96 		64'h5bd82ab37fd3d86c
`define	S97 		64'he4a057e7dba678f8
`define	S98 		64'ha940ed4eb768b951
`define	S99 		64'h73811a9d4af1fba3
`define	S100 		64'h940337bb95c23ce6
`define	S101 		64'h38076df62f84756d
`define	S102 		64'h400f9b6c7b0caffa
`define	S103 		64'hc01eb4d8d61dd054
`define	S104 		64'hc02de931a83e60a9
`define	S105 		64'hc05a1262705881f3
`define	S106 		64'hc0a426c4c0b18247
`define	S107 		64'hc1484f098142868f
`define	S108 		64'hc390dc1202858b9f
`define	S109 		64'hc4317824050e9cbf
`define	S110 		64'hc873b0480e19b5df
`define	S111 		64'hd0f6e0901832ee3f
`define	S112 		64'hf1fd01a03045125f
`define	S113 		64'h92eb03c0408f26bf
`define	S114 		64'h37d70500811b4bdf
`define	S115 		64'h5cbf0a010237dc3e
`define	S116 		64'he96f1603044a745c
`define	S117 		64'hb3df2e070c94acb9
`define	S118 		64'h54af5e0f1d2dd5d3
`define	S119 		64'hf95ffe1f3e7e6e26
`define	S120 		64'h83ae3e3f58d8926d
`define	S121 		64'h045c7e7fb1b1a6fb
`define	S122 		64'h08a8befe4342cb56
`define	S123 		64'h1151ff7c86855dac
`define	S124 		64'h33b23cf9090ff6f8
`define	S125 		64'h54747973121a2b50
`define	S126 		64'hf8f8b2e724345da0
`define	S127 		64'h81e1e74f6c4cf6e1
`define	S128 		64'h02c20c9ffc9d2b63
`define	S129 		64'h078419bedd3f5de6
`define	S130 		64'h0c0833fdbe5bf66c
`define	S131 		64'h1810657a58b62af8
`define	S132 		64'h20308af4b1485f50
`define	S133 		64'h607197694290f1a0
`define	S134 		64'ha0f2acd3852122e0
`define	S135 		64'h61f5d9260e634761
`define	S136 		64'ha2fa724c18e7c9e2
`define	S137 		64'h67e4a69831ea5a65
`define	S138 		64'hacc9cfb043f4feea
`define	S139		64'h79925de087cd3375
`define	S140 		64'h8234fb410b9f65ca
`define	S141 		64'h06793483173b8e15
`define	S142 		64'h0ee369872a56922a
`define	S143 		64'h1fc7938f74a9a674
`define	S144 		64'h2c8ea59fcd72cac8
`define	S145 		64'h791dcbbe9ec55f10
`define	S146 		64'h832a55fd398ff120
`define	S147 		64'h0554eb7b531a2361
`define	S148 		64'h0bb914f7a63445e2
`define	S149 		64'h1463296e684cce64
`define	S150 		64'h38c752dcf09d52e8
`define	S151 		64'h418fe739c13fe770
`define	S152 		64'hc21e0c72825a09c0
`define	S153 		64'hc62c18e504b41a01
`define	S154 		64'hce58314b0d4c3e03
`define	S155 		64'hdea062971e9c7207
`define	S156 		64'hef4087af393ca60f
`define	S157 		64'hbd818ddf525dca1f
`define	S158 		64'h4a029b3fa4be5e3f
`define	S159 		64'hd605b47e6d58f25e
`define	S160 		64'hfe0ae8fcfeb126bd
`define	S161 		64'h8e151179d9434bdb
`define	S162 		64'h1e3b22f2b287dc37
`define	S163 		64'h2e674765450a744e
`define	S164 		64'h7ecfcccb8e14ac9c
`define	S165 		64'h8f9e5916182dd5b8
`define	S166 		64'h1c2cf22c307e6ed1
`define	S167 		64'h2859265840d89322

//S_array[168*w-1:0] 
`define S_array     {`S167,`S166,`S165,`S164,`S163,`S162,`S161,`S160,`S159,`S158,`S157,`S156,`S155,`S154,`S153,`S152,`S151,`S150,`S149,`S148,`S147,`S146,`S145,`S144,`S143,`S142,`S141,`S140,`S139,`S138,`S137,`S136,`S135,`S134,`S133,`S132,`S131,`S130,`S129,`S128,`S127,`S126,`S125,`S124,`S123,`S122,`S121,`S120,`S119,`S118,`S117,`S116,`S115,`S114,`S113,`S112,`S111,`S110,`S109,`S108,`S107,`S106,`S105,`S104,`S103,`S102,`S101,`S100,`S99 ,`S98 , `S97 ,`S96 ,`S95 ,`S94 ,`S93 ,`S92 ,`S91 ,`S90 ,`S89 ,`S88 ,`S87 ,`S86 ,`S85 ,`S84 ,`S83 ,`S82 ,`S81 ,`S80 ,`S79 ,`S78 ,`S77 ,`S76 ,`S75 ,`S74 ,`S73 ,`S72 ,`S71 ,`S70 , `S69 ,`S68 ,`S67 ,`S66 ,`S65 ,`S64 ,`S63 ,`S62 ,`S61 ,`S60 ,`S59 ,`S58 ,`S57 ,`S56 ,`S55 ,`S54 ,`S53 ,`S52 ,`S51 ,`S50 ,`S49 ,`S48 ,`S47 ,`S46 ,`S45 ,`S44 ,`S43 ,`S42 ,`S41 ,`S40 ,`S39 ,`S38 ,`S37 ,`S36 ,`S35 ,`S34 ,`S33 ,`S32 ,`S31 ,`S30 ,`S29 ,`S28 ,`S27 ,`S26 ,`S25 ,`S24 ,`S23 ,`S22 ,`S21 ,`S20 ,`S19 ,`S18 ,`S17 ,`S16 ,`S15 ,`S14 ,`S13 ,`S12 ,`S11 ,`S10 ,`S9  ,`S8  ,`S7  ,`S6  ,`S5  ,`S4  ,`S3  ,`S2  ,`S1  ,`S0  }
//t
`define t0	8'd17
`define t1	8'd18
`define t2	8'd21
`define t3	8'd31
`define t4	8'd67
//t_array[5*byte-1:0]
`define t_array     {`t0,`t1,`t2,`t3,`t4}

//shift amounts
//r(i-n)
`define r0		8'd10
`define r1		8'd5
`define r2		8'd13
`define r3		8'd10
`define r4		8'd11
`define r5		8'd12
`define r6		8'd2
`define r7		8'd7
`define r8		8'd14
`define r9		8'd15
`define r10		8'd7
`define r11		8'd13
`define r12		8'd11
`define r13		8'd7
`define r14		8'd6
`define r15		8'd12

//r_array[16*byte-1:0]
`define r_array     {`r15,`r14,`r13,`r12,`r11,`r10,`r9,`r8,`r7,`r6,`r5,`r4,`r3,`r2,`r1,`r0}

//l(i-n)
`define l0		8'd11
`define l1		8'd24
`define l2		8'd9
`define l3		8'd16
`define l4		8'd15
`define l5		8'd9
`define l6		8'd27
`define l7		8'd15
`define l8		8'd6
`define l9		8'd2
`define l10		8'd29
`define l11		8'd8
`define l12		8'd15
`define l13		8'd5
`define l14		8'd31
`define l15		8'd9

//l_array[16*byte-1:0]
`define l_array     {`l15,`l14,`l13,`l12,`l11,`l10,`l9,`l8,`l7,`l6,`l5,`l4,`l3,`l2,`l1,`l0}

`define clog2(x)\
(x == 0) ? 0   : (x<16**1) ? 4: (x<16**2) ? 8: (x<16**3) ? 12: (x<16**4) ? 16: (x<16**5) ? 20: (x<16**6) ? 24: (x<16**7) ? 28: (x<16**8) ? 32: (x<16**9) ? 36: (x<16**10) ? 40: (x<16**11) ? 44: (x<16**12) ? 48: (x<16**13) ? 52: (x<16**14) ? 56: (x<16**15) ? 60: (x<16**16) ? 64: (x<16**17) ? 68: (x<16**18) ? 72: (x<16**19) ? 76: (x<16**20) ? 80: (x<16**21) ? 84: (x<16**22) ? 88: (x<16**23) ? 92: (x<16**24) ? 96: (x<16**25) ? 100: (x<16**26) ? 104: (x<16**27) ? 108: (x<16**28) ? 112: (x<16**29) ? 116: (x<16**30) ? 120: (x<16**31) ? 124: (x<16**32) ? 128: (x<16**33) ? 132: (x<16**34) ? 136: (x<16**35) ? 140: (x<16**36) ? 144: (x<16**37) ? 148: (x<16**38) ? 152: (x<16**39) ? 156: (x<16**40) ? 160: (x<16**41) ? 164: (x<16**42) ? 168: (x<16**43) ? 172: (x<16**44) ? 176: (x<16**45) ? 180: (x<16**46) ? 184: (x<16**47) ? 188: (x<16**48) ? 192: (x<16**49) ? 196: (x<16**50) ? 200: (x<16**51) ? 204: (x<16**52) ? 208: (x<16**53) ? 212: (x<16**54) ? 216: (x<16**55) ? 220: (x<16**56) ? 224: (x<16**57) ? 228: (x<16**58) ? 232: (x<16**59) ? 236: (x<16**60) ? 240: (x<16**61) ? 244: (x<16**62) ? 248: (x<16**63) ? 252: (x<16**64) ? 256: (x<16**65) ? 260: (x<16**66) ? 264: (x<16**67) ? 268: (x<16**68) ? 272: (x<16**69) ? 276: (x<16**70) ? 280: (x<16**71) ? 284: (x<16**72) ? 288: (x<16**73) ? 292: (x<16**74) ? 296: (x<16**75) ? 300: (x<16**76) ? 304: (x<16**77) ? 308: (x<16**78) ? 312: (x<16**79) ? 316: (x<16**80) ? 320: (x<16**81) ? 324: (x<16**82) ? 328: (x<16**83) ? 332: (x<16**84) ? 336: (x<16**85) ? 340: (x<16**86) ? 344: (x<16**87) ? 348: (x<16**88) ? 352: (x<16**89) ? 356: (x<16**90) ? 360: (x<16**91) ? 364: (x<16**92) ? 368: (x<16**93) ? 372: (x<16**94) ? 376: (x<16**95) ? 380: (x<16**96) ? 384: (x<16**97) ? 388: (x<16**98) ? 392: (x<16**99) ? 396: (x<16**100) ? 400: (x<16**101) ? 404: (x<16**102) ? 408: (x<16**103) ? 412: (x<16**104) ? 416: (x<16**105) ? 420: (x<16**106) ? 424: (x<16**107) ? 428: (x<16**108) ? 432: (x<16**109) ? 436: (x<16**110) ? 440: (x<16**111) ? 444: (x<16**112) ? 448: (x<16**113) ? 452: (x<16**114) ? 456: (x<16**115) ? 460: (x<16**116) ? 464: (x<16**117) ? 468: (x<16**118) ? 472: (x<16**119) ? 476: (x<16**120) ? 480: (x<16**121) ? 484: (x<16**122) ? 488: (x<16**123) ? 492: (x<16**124) ? 496: (x<16**125) ? 500: (x<16**126) ? 504: (x<16**127) ? 508: (x<16**128) ? 512: (x<16**129) ? 516: (x<16**130) ? 520: (x<16**131) ? 524: (x<16**132) ? 528: (x<16**133) ? 532: (x<16**134) ? 536: (x<16**135) ? 540: (x<16**136) ? 544: (x<16**137) ? 548: (x<16**138) ? 552: (x<16**139) ? 556: (x<16**140) ? 560: (x<16**141) ? 564: (x<16**142) ? 568: (x<16**143) ? 572: (x<16**144) ? 576: (x<16**145) ? 580: (x<16**146) ? 584: (x<16**147) ? 588: (x<16**148) ? 592: (x<16**149) ? 596: (x<16**150) ? 600: (x<16**151) ? 604: (x<16**152) ? 608: (x<16**153) ? 612: (x<16**154) ? 616: (x<16**155) ? 620: (x<16**156) ? 624: (x<16**157) ? 628: (x<16**158) ? 632: (x<16**159) ? 636: (x<16**160) ? 640: (x<16**161) ? 644: (x<16**162) ? 648: (x<16**163) ? 652: (x<16**164) ? 656: (x<16**165) ? 660: (x<16**166) ? 664: (x<16**167) ? 668: (x<16**168) ? 672: (x<16**169) ? 676: (x<16**170) ? 680: (x<16**171) ? 684: (x<16**172) ? 688: (x<16**173) ? 692: (x<16**174) ? 696: (x<16**175) ? 700: (x<16**176) ? 704: (x<16**177) ? 708: (x<16**178) ? 712: (x<16**179) ? 716: (x<16**180) ? 720: (x<16**181) ? 724: (x<16**182) ? 728: (x<16**183) ? 732: (x<16**184) ? 736: (x<16**185) ? 740: (x<16**186) ? 744: (x<16**187) ? 748: (x<16**188) ? 752: (x<16**189) ? 756: (x<16**190) ? 760: (x<16**191) ? 764: (x<16**192) ? 768: (x<16**193) ? 772: (x<16**194) ? 776: (x<16**195) ? 780: (x<16**196) ? 784: (x<16**197) ? 788: (x<16**198) ? 792: (x<16**199) ? 796: (x<16**200) ? 800: (x<16**201) ? 804: (x<16**202) ? 808: (x<16**203) ? 812: (x<16**204) ? 816: (x<16**205) ? 820: (x<16**206) ? 824: (x<16**207) ? 828: (x<16**208) ? 832: (x<16**209) ? 836: (x<16**210) ? 840: (x<16**211) ? 844: (x<16**212) ? 848: (x<16**213) ? 852: (x<16**214) ? 856: (x<16**215) ? 860: (x<16**216) ? 864: (x<16**217) ? 868: (x<16**218) ? 872: (x<16**219) ? 876: (x<16**220) ? 880: (x<16**221) ? 884: (x<16**222) ? 888: (x<16**223) ? 892: (x<16**224) ? 896: (x<16**225) ? 900: (x<16**226) ? 904: (x<16**227) ? 908: (x<16**228) ? 912: (x<16**229) ? 916: (x<16**230) ? 920: (x<16**231) ? 924: (x<16**232) ? 928: (x<16**233) ? 932: (x<16**234) ? 936: (x<16**235) ? 940: (x<16**236) ? 944: (x<16**237) ? 948: (x<16**238) ? 952: (x<16**239) ? 956: (x<16**240) ? 960: (x<16**241) ? 964: (x<16**242) ? 968: (x<16**243) ? 972: (x<16**244) ? 976: (x<16**245) ? 980: (x<16**246) ? 984: (x<16**247) ? 988: (x<16**248) ? 992: (x<16**249) ? 996: (x<16**250) ? 1000: (x<16**251) ? 1004: (x<16**252) ? 1008: (x<16**253) ? 1012: (x<16**254) ? 1016: (x<16**255) ? 1020: (x<16**256) ? 1024: (x<16**257) ? 1028: (x<16**258) ? 1032: (x<16**259) ? 1036: (x<16**260) ? 1040: (x<16**261) ? 1044: (x<16**262) ? 1048: (x<16**263) ? 1052: (x<16**264) ? 1056: (x<16**265) ? 1060: (x<16**266) ? 1064: (x<16**267) ? 1068: (x<16**268) ? 1072: (x<16**269) ? 1076: (x<16**270) ? 1080: (x<16**271) ? 1084: (x<16**272) ? 1088: (x<16**273) ? 1092: (x<16**274) ? 1096: (x<16**275) ? 1100: (x<16**276) ? 1104: (x<16**277) ? 1108: (x<16**278) ? 1112: (x<16**279) ? 1116: (x<16**280) ? 1120: (x<16**281) ? 1124: (x<16**282) ? 1128: (x<16**283) ? 1132: (x<16**284) ? 1136: (x<16**285) ? 1140: (x<16**286) ? 1144: (x<16**287) ? 1148: (x<16**288) ? 1152: (x<16**289) ? 1156: (x<16**290) ? 1160: (x<16**291) ? 1164: (x<16**292) ? 1168: (x<16**293) ? 1172: (x<16**294) ? 1176: (x<16**295) ? 1180: (x<16**296) ? 1184: (x<16**297) ? 1188: (x<16**298) ? 1192: (x<16**299) ? 1196: (x<16**300) ? 1200: (x<16**301) ? 1204: (x<16**302) ? 1208: (x<16**303) ? 1212: (x<16**304) ? 1216: (x<16**305) ? 1220: (x<16**306) ? 1224: (x<16**307) ? 1228: (x<16**308) ? 1232: (x<16**309) ? 1236: (x<16**310) ? 1240: (x<16**311) ? 1244: (x<16**312) ? 1248: (x<16**313) ? 1252: (x<16**314) ? 1256: (x<16**315) ? 1260: (x<16**316) ? 1264: (x<16**317) ? 1268: (x<16**318) ? 1272: (x<16**319) ? 1276: (x<16**320) ? 1280: (x<16**321) ? 1284: (x<16**322) ? 1288: (x<16**323) ? 1292: (x<16**324) ? 1296: (x<16**325) ? 1300: (x<16**326) ? 1304: (x<16**327) ? 1308: (x<16**328) ? 1312: (x<16**329) ? 1316: (x<16**330) ? 1320: (x<16**331) ? 1324: (x<16**332) ? 1328: (x<16**333) ? 1332: (x<16**334) ? 1336: (x<16**335) ? 1340: (x<16**336) ? 1344: (x<16**337) ? 1348: (x<16**338) ? 1352: (x<16**339) ? 1356: (x<16**340) ? 1360: (x<16**341) ? 1364: (x<16**342) ? 1368: (x<16**343) ? 1372: (x<16**344) ? 1376: (x<16**345) ? 1380: (x<16**346) ? 1384: (x<16**347) ? 1388: (x<16**348) ? 1392: (x<16**349) ? 1396: (x<16**350) ? 1400: (x<16**351) ? 1404: (x<16**352) ? 1408: (x<16**353) ? 1412: (x<16**354) ? 1416: (x<16**355) ? 1420: (x<16**356) ? 1424: (x<16**357) ? 1428: (x<16**358) ? 1432: (x<16**359) ? 1436: (x<16**360) ? 1440: (x<16**361) ? 1444: (x<16**362) ? 1448: (x<16**363) ? 1452: (x<16**364) ? 1456: (x<16**365) ? 1460: (x<16**366) ? 1464: (x<16**367) ? 1468: (x<16**368) ? 1472: (x<16**369) ? 1476: (x<16**370) ? 1480: (x<16**371) ? 1484: (x<16**372) ? 1488: (x<16**373) ? 1492: (x<16**374) ? 1496: (x<16**375) ? 1500: (x<16**376) ? 1504: (x<16**377) ? 1508: (x<16**378) ? 1512: (x<16**379) ? 1516: (x<16**380) ? 1520: (x<16**381) ? 1524: (x<16**382) ? 1528: (x<16**383) ? 1532: (x<16**384) ? 1536: (x<16**385) ? 1540: (x<16**386) ? 1544: (x<16**387) ? 1548: (x<16**388) ? 1552: (x<16**389) ? 1556: (x<16**390) ? 1560: (x<16**391) ? 1564: (x<16**392) ? 1568: (x<16**393) ? 1572: (x<16**394) ? 1576: (x<16**395) ? 1580: (x<16**396) ? 1584: (x<16**397) ? 1588: (x<16**398) ? 1592: (x<16**399) ? 1596: (x<16**400) ? 1600: (x<16**401) ? 1604: (x<16**402) ? 1608: (x<16**403) ? 1612: (x<16**404) ? 1616: (x<16**405) ? 1620: (x<16**406) ? 1624: (x<16**407) ? 1628: (x<16**408) ? 1632: (x<16**409) ? 1636: (x<16**410) ? 1640: (x<16**411) ? 1644: (x<16**412) ? 1648: (x<16**413) ? 1652: (x<16**414) ? 1656: (x<16**415) ? 1660: (x<16**416) ? 1664: (x<16**417) ? 1668: (x<16**418) ? 1672: (x<16**419) ? 1676: (x<16**420) ? 1680: (x<16**421) ? 1684: (x<16**422) ? 1688: (x<16**423) ? 1692: (x<16**424) ? 1696: (x<16**425) ? 1700: (x<16**426) ? 1704: (x<16**427) ? 1708: (x<16**428) ? 1712: (x<16**429) ? 1716: (x<16**430) ? 1720: (x<16**431) ? 1724: (x<16**432) ? 1728: (x<16**433) ? 1732: (x<16**434) ? 1736: (x<16**435) ? 1740: (x<16**436) ? 1744: (x<16**437) ? 1748: (x<16**438) ? 1752: (x<16**439) ? 1756: (x<16**440) ? 1760: (x<16**441) ? 1764: (x<16**442) ? 1768: (x<16**443) ? 1772: (x<16**444) ? 1776: (x<16**445) ? 1780: (x<16**446) ? 1784: (x<16**447) ? 1788: (x<16**448) ? 1792: (x<16**449) ? 1796: (x<16**450) ? 1800: (x<16**451) ? 1804: (x<16**452) ? 1808: (x<16**453) ? 1812: (x<16**454) ? 1816: (x<16**455) ? 1820: (x<16**456) ? 1824: (x<16**457) ? 1828: (x<16**458) ? 1832: (x<16**459) ? 1836: (x<16**460) ? 1840: (x<16**461) ? 1844: (x<16**462) ? 1848: (x<16**463) ? 1852: (x<16**464) ? 1856: (x<16**465) ? 1860: (x<16**466) ? 1864: (x<16**467) ? 1868: (x<16**468) ? 1872: (x<16**469) ? 1876: (x<16**470) ? 1880: (x<16**471) ? 1884: (x<16**472) ? 1888: (x<16**473) ? 1892: (x<16**474) ? 1896: (x<16**475) ? 1900: (x<16**476) ? 1904: (x<16**477) ? 1908: (x<16**478) ? 1912: (x<16**479) ? 1916: (x<16**480) ? 1920: (x<16**481) ? 1924: (x<16**482) ? 1928: (x<16**483) ? 1932: (x<16**484) ? 1936: (x<16**485) ? 1940: (x<16**486) ? 1944: (x<16**487) ? 1948: (x<16**488) ? 1952: (x<16**489) ? 1956: (x<16**490) ? 1960: (x<16**491) ? 1964: (x<16**492) ? 1968: (x<16**493) ? 1972: (x<16**494) ? 1976: (x<16**495) ? 1980: (x<16**496) ? 1984: (x<16**497) ? 1988: (x<16**498) ? 1992: (x<16**499) ? 1996: (x<16**500) ? 2000: (x<16**501) ? 2004: (x<16**502) ? 2008: (x<16**503) ? 2012: (x<16**504) ? 2016: (x<16**505) ? 2020: (x<16**506) ? 2024: (x<16**507) ? 2028: (x<16**508) ? 2032: (x<16**509) ? 2036: (x<16**510) ? 2040: (x<16**511) ? 2044: (x<16**512) ? 2048: (x<16**513) ? 2052: (x<16**514) ? 2056: (x<16**515) ? 2060: (x<16**516) ? 2064: (x<16**517) ? 2068: (x<16**518) ? 2072: (x<16**519) ? 2076: (x<16**520) ? 2080: (x<16**521) ? 2084: (x<16**522) ? 2088: (x<16**523) ? 2092: (x<16**524) ? 2096: (x<16**525) ? 2100: (x<16**526) ? 2104: (x<16**527) ? 2108: (x<16**528) ? 2112: (x<16**529) ? 2116: (x<16**530) ? 2120: (x<16**531) ? 2124: (x<16**532) ? 2128: (x<16**533) ? 2132: (x<16**534) ? 2136: (x<16**535) ? 2140: (x<16**536) ? 2144: (x<16**537) ? 2148: (x<16**538) ? 2152: (x<16**539) ? 2156: (x<16**540) ? 2160: (x<16**541) ? 2164: (x<16**542) ? 2168: (x<16**543) ? 2172: (x<16**544) ? 2176: (x<16**545) ? 2180: (x<16**546) ? 2184: (x<16**547) ? 2188: (x<16**548) ? 2192: (x<16**549) ? 2196: (x<16**550) ? 2200: (x<16**551) ? 2204: (x<16**552) ? 2208: (x<16**553) ? 2212: (x<16**554) ? 2216: (x<16**555) ? 2220: (x<16**556) ? 2224: (x<16**557) ? 2228: (x<16**558) ? 2232: (x<16**559) ? 2236: (x<16**560) ? 2240: (x<16**561) ? 2244: (x<16**562) ? 2248: (x<16**563) ? 2252: (x<16**564) ? 2256: (x<16**565) ? 2260: (x<16**566) ? 2264: (x<16**567) ? 2268: (x<16**568) ? 2272: (x<16**569) ? 2276: (x<16**570) ? 2280: (x<16**571) ? 2284: (x<16**572) ? 2288: (x<16**573) ? 2292: (x<16**574) ? 2296: (x<16**575) ? 2300: (x<16**576) ? 2304: (x<16**577) ? 2308: (x<16**578) ? 2312: (x<16**579) ? 2316: (x<16**580) ? 2320: (x<16**581) ? 2324: (x<16**582) ? 2328: (x<16**583) ? 2332: (x<16**584) ? 2336: (x<16**585) ? 2340: (x<16**586) ? 2344: (x<16**587) ? 2348: (x<16**588) ? 2352: (x<16**589) ? 2356: (x<16**590) ? 2360: (x<16**591) ? 2364: (x<16**592) ? 2368: (x<16**593) ? 2372: (x<16**594) ? 2376: (x<16**595) ? 2380: (x<16**596) ? 2384: (x<16**597) ? 2388: (x<16**598) ? 2392: (x<16**599) ? 2396: (x<16**600) ? 2400: (x<16**601) ? 2404: (x<16**602) ? 2408: (x<16**603) ? 2412: (x<16**604) ? 2416: (x<16**605) ? 2420: (x<16**606) ? 2424: (x<16**607) ? 2428: (x<16**608) ? 2432: (x<16**609) ? 2436: (x<16**610) ? 2440: (x<16**611) ? 2444: (x<16**612) ? 2448: (x<16**613) ? 2452: (x<16**614) ? 2456: (x<16**615) ? 2460: (x<16**616) ? 2464: (x<16**617) ? 2468: (x<16**618) ? 2472: (x<16**619) ? 2476: (x<16**620) ? 2480: (x<16**621) ? 2484: (x<16**622) ? 2488: (x<16**623) ? 2492: (x<16**624) ? 2496: (x<16**625) ? 2500: (x<16**626) ? 2504: (x<16**627) ? 2508: (x<16**628) ? 2512: (x<16**629) ? 2516: (x<16**630) ? 2520: (x<16**631) ? 2524: (x<16**632) ? 2528: (x<16**633) ? 2532: (x<16**634) ? 2536: (x<16**635) ? 2540: (x<16**636) ? 2544: (x<16**637) ? 2548: (x<16**638) ? 2552: (x<16**639) ? 2556: (x<16**640) ? 2560: (x<16**641) ? 2564: (x<16**642) ? 2568: (x<16**643) ? 2572: (x<16**644) ? 2576: (x<16**645) ? 2580: (x<16**646) ? 2584: (x<16**647) ? 2588: (x<16**648) ? 2592: (x<16**649) ? 2596: (x<16**650) ? 2600: (x<16**651) ? 2604: (x<16**652) ? 2608: (x<16**653) ? 2612: (x<16**654) ? 2616: (x<16**655) ? 2620: (x<16**656) ? 2624: (x<16**657) ? 2628: (x<16**658) ? 2632: (x<16**659) ? 2636: (x<16**660) ? 2640: (x<16**661) ? 2644: (x<16**662) ? 2648: (x<16**663) ? 2652: (x<16**664) ? 2656: (x<16**665) ? 2660: (x<16**666) ? 2664: (x<16**667) ? 2668: (x<16**668) ? 2672: (x<16**669) ? 2676: (x<16**670) ? 2680: (x<16**671) ? 2684: (x<16**672) ? 2688: (x<16**673) ? 2692: (x<16**674) ? 2696: (x<16**675) ? 2700: (x<16**676) ? 2704: (x<16**677) ? 2708: (x<16**678) ? 2712: (x<16**679) ? 2716: (x<16**680) ? 2720: (x<16**681) ? 2724: (x<16**682) ? 2728: (x<16**683) ? 2732: (x<16**684) ? 2736: (x<16**685) ? 2740: (x<16**686) ? 2744: (x<16**687) ? 2748: (x<16**688) ? 2752: (x<16**689) ? 2756: (x<16**690) ? 2760: (x<16**691) ? 2764: (x<16**692) ? 2768: (x<16**693) ? 2772: (x<16**694) ? 2776: (x<16**695) ? 2780: (x<16**696) ? 2784: (x<16**697) ? 2788: (x<16**698) ? 2792: (x<16**699) ? 2796: (x<16**700) ? 2800: (x<16**701) ? 2804: (x<16**702) ? 2808: (x<16**703) ? 2812: (x<16**704) ? 2816: (x<16**705) ? 2820: (x<16**706) ? 2824: (x<16**707) ? 2828: (x<16**708) ? 2832: (x<16**709) ? 2836: (x<16**710) ? 2840: (x<16**711) ? 2844: (x<16**712) ? 2848: (x<16**713) ? 2852: (x<16**714) ? 2856: (x<16**715) ? 2860: (x<16**716) ? 2864: (x<16**717) ? 2868: (x<16**718) ? 2872: (x<16**719) ? 2876: (x<16**720) ? 2880: (x<16**721) ? 2884: (x<16**722) ? 2888: (x<16**723) ? 2892: (x<16**724) ? 2896: (x<16**725) ? 2900: (x<16**726) ? 2904: (x<16**727) ? 2908: (x<16**728) ? 2912: (x<16**729) ? 2916: (x<16**730) ? 2920: (x<16**731) ? 2924: (x<16**732) ? 2928: (x<16**733) ? 2932: (x<16**734) ? 2936: (x<16**735) ? 2940: (x<16**736) ? 2944: (x<16**737) ? 2948: (x<16**738) ? 2952: (x<16**739) ? 2956: (x<16**740) ? 2960: (x<16**741) ? 2964: (x<16**742) ? 2968: (x<16**743) ? 2972: (x<16**744) ? 2976: (x<16**745) ? 2980: (x<16**746) ? 2984: (x<16**747) ? 2988: (x<16**748) ? 2992: (x<16**749) ? 2996: (x<16**750) ? 3000: (x<16**751) ? 3004: (x<16**752) ? 3008: (x<16**753) ? 3012: (x<16**754) ? 3016: (x<16**755) ? 3020: (x<16**756) ? 3024: (x<16**757) ? 3028: (x<16**758) ? 3032: (x<16**759) ? 3036: (x<16**760) ? 3040: (x<16**761) ? 3044: (x<16**762) ? 3048: (x<16**763) ? 3052: (x<16**764) ? 3056: (x<16**765) ? 3060: (x<16**766) ? 3064: (x<16**767) ? 3068: (x<16**768) ? 3072: (x<16**769) ? 3076: (x<16**770) ? 3080: (x<16**771) ? 3084: (x<16**772) ? 3088: (x<16**773) ? 3092: (x<16**774) ? 3096: (x<16**775) ? 3100: (x<16**776) ? 3104: (x<16**777) ? 3108: (x<16**778) ? 3112: (x<16**779) ? 3116: (x<16**780) ? 3120: (x<16**781) ? 3124: (x<16**782) ? 3128: (x<16**783) ? 3132: (x<16**784) ? 3136: (x<16**785) ? 3140: (x<16**786) ? 3144: (x<16**787) ? 3148: (x<16**788) ? 3152: (x<16**789) ? 3156: (x<16**790) ? 3160: (x<16**791) ? 3164: (x<16**792) ? 3168: (x<16**793) ? 3172: (x<16**794) ? 3176: (x<16**795) ? 3180: (x<16**796) ? 3184: (x<16**797) ? 3188: (x<16**798) ? 3192: (x<16**799) ? 3196: (x<16**800) ? 3200: (x<16**801) ? 3204: (x<16**802) ? 3208: (x<16**803) ? 3212: (x<16**804) ? 3216: (x<16**805) ? 3220: (x<16**806) ? 3224: (x<16**807) ? 3228: (x<16**808) ? 3232: (x<16**809) ? 3236: (x<16**810) ? 3240: (x<16**811) ? 3244: (x<16**812) ? 3248: (x<16**813) ? 3252: (x<16**814) ? 3256: (x<16**815) ? 3260: (x<16**816) ? 3264: (x<16**817) ? 3268: (x<16**818) ? 3272: (x<16**819) ? 3276: (x<16**820) ? 3280: (x<16**821) ? 3284: (x<16**822) ? 3288: (x<16**823) ? 3292: (x<16**824) ? 3296: (x<16**825) ? 3300: (x<16**826) ? 3304: (x<16**827) ? 3308: (x<16**828) ? 3312: (x<16**829) ? 3316: (x<16**830) ? 3320: (x<16**831) ? 3324: (x<16**832) ? 3328: (x<16**833) ? 3332: (x<16**834) ? 3336: (x<16**835) ? 3340: (x<16**836) ? 3344: (x<16**837) ? 3348: (x<16**838) ? 3352: (x<16**839) ? 3356: (x<16**840) ? 3360: (x<16**841) ? 3364: (x<16**842) ? 3368: (x<16**843) ? 3372: (x<16**844) ? 3376: (x<16**845) ? 3380: (x<16**846) ? 3384: (x<16**847) ? 3388: (x<16**848) ? 3392: (x<16**849) ? 3396: (x<16**850) ? 3400: (x<16**851) ? 3404: (x<16**852) ? 3408: (x<16**853) ? 3412: (x<16**854) ? 3416: (x<16**855) ? 3420: (x<16**856) ? 3424: (x<16**857) ? 3428: (x<16**858) ? 3432: (x<16**859) ? 3436: (x<16**860) ? 3440: (x<16**861) ? 3444: (x<16**862) ? 3448: (x<16**863) ? 3452: (x<16**864) ? 3456: (x<16**865) ? 3460: (x<16**866) ? 3464: (x<16**867) ? 3468: (x<16**868) ? 3472: (x<16**869) ? 3476: (x<16**870) ? 3480: (x<16**871) ? 3484: (x<16**872) ? 3488: (x<16**873) ? 3492: (x<16**874) ? 3496: (x<16**875) ? 3500: (x<16**876) ? 3504: (x<16**877) ? 3508: (x<16**878) ? 3512: (x<16**879) ? 3516: (x<16**880) ? 3520: (x<16**881) ? 3524: (x<16**882) ? 3528: (x<16**883) ? 3532: (x<16**884) ? 3536: (x<16**885) ? 3540: (x<16**886) ? 3544: (x<16**887) ? 3548: (x<16**888) ? 3552: (x<16**889) ? 3556: (x<16**890) ? 3560: (x<16**891) ? 3564: (x<16**892) ? 3568: (x<16**893) ? 3572: (x<16**894) ? 3576: (x<16**895) ? 3580: (x<16**896) ? 3584: (x<16**897) ? 3588: (x<16**898) ? 3592: (x<16**899) ? 3596: (x<16**900) ? 3600: (x<16**901) ? 3604: (x<16**902) ? 3608: (x<16**903) ? 3612: (x<16**904) ? 3616: (x<16**905) ? 3620: (x<16**906) ? 3624: (x<16**907) ? 3628: (x<16**908) ? 3632: (x<16**909) ? 3636: (x<16**910) ? 3640: (x<16**911) ? 3644: (x<16**912) ? 3648: (x<16**913) ? 3652: (x<16**914) ? 3656: (x<16**915) ? 3660: (x<16**916) ? 3664: (x<16**917) ? 3668: (x<16**918) ? 3672: (x<16**919) ? 3676: (x<16**920) ? 3680: (x<16**921) ? 3684: (x<16**922) ? 3688: (x<16**923) ? 3692: (x<16**924) ? 3696: (x<16**925) ? 3700: (x<16**926) ? 3704: (x<16**927) ? 3708: (x<16**928) ? 3712: (x<16**929) ? 3716: (x<16**930) ? 3720: (x<16**931) ? 3724: (x<16**932) ? 3728: (x<16**933) ? 3732: (x<16**934) ? 3736: (x<16**935) ? 3740: (x<16**936) ? 3744: (x<16**937) ? 3748: (x<16**938) ? 3752: (x<16**939) ? 3756: (x<16**940) ? 3760: (x<16**941) ? 3764: (x<16**942) ? 3768: (x<16**943) ? 3772: (x<16**944) ? 3776: (x<16**945) ? 3780: (x<16**946) ? 3784: (x<16**947) ? 3788: (x<16**948) ? 3792: (x<16**949) ? 3796: (x<16**950) ? 3800: (x<16**951) ? 3804: (x<16**952) ? 3808: (x<16**953) ? 3812: (x<16**954) ? 3816: (x<16**955) ? 3820: (x<16**956) ? 3824: (x<16**957) ? 3828: (x<16**958) ? 3832: (x<16**959) ? 3836: (x<16**960) ? 3840: (x<16**961) ? 3844: (x<16**962) ? 3848: (x<16**963) ? 3852: (x<16**964) ? 3856: (x<16**965) ? 3860: (x<16**966) ? 3864: (x<16**967) ? 3868: (x<16**968) ? 3872: (x<16**969) ? 3876: (x<16**970) ? 3880: (x<16**971) ? 3884: (x<16**972) ? 3888: (x<16**973) ? 3892: (x<16**974) ? 3896: (x<16**975) ? 3900: (x<16**976) ? 3904: (x<16**977) ? 3908: (x<16**978) ? 3912: (x<16**979) ? 3916: (x<16**980) ? 3920: (x<16**981) ? 3924: (x<16**982) ? 3928: (x<16**983) ? 3932: (x<16**984) ? 3936: (x<16**985) ? 3940: (x<16**986) ? 3944: (x<16**987) ? 3948: (x<16**988) ? 3952: (x<16**989) ? 3956: (x<16**990) ? 3960: (x<16**991) ? 3964: (x<16**992) ? 3968: (x<16**993) ? 3972: (x<16**994) ? 3976: (x<16**995) ? 3980: (x<16**996) ? 3984: (x<16**997) ? 3988: (x<16**998) ? 3992: (x<16**999) ? 3996: (x<16**1000) ? 4000: (x<16**1001) ? 4004: (x<16**1002) ? 4008: (x<16**1003) ? 4012: (x<16**1004) ? 4016: (x<16**1005) ? 4020: (x<16**1006) ? 4024: (x<16**1007) ? 4028: (x<16**1008) ? 4032: (x<16**1009) ? 4036: (x<16**1010) ? 4040: (x<16**1011) ? 4044: (x<16**1012) ? 4048: (x<16**1013) ? 4052: (x<16**1014) ? 4056: (x<16**1015) ? 4060: (x<16**1016) ? 4064: (x<16**1017) ? 4068: (x<16**1018) ? 4072: (x<16**1019) ? 4076: (x<16**1020) ? 4080: (x<16**1021) ? 4084: (x<16**1022) ? 4088: (x<16**1023) ? 4092: (x<16**1024) ? 4096 : -1



`define padding(x)\
(x == 0) ? 4096 : (x < 16**1) ? 4092 : (x < 16**2) ? 4088 : (x < 16**3) ? 4084 : (x < 16**4) ? 4080 : (x < 16**5) ? 4076 : (x < 16**6) ? 4072 : (x < 16**7) ? 4068 : (x < 16**8) ? 4064 : (x < 16**9) ? 4060 : (x < 16**10) ? 4056 : (x < 16**11) ? 4052 : (x < 16**12) ? 4048 : (x < 16**13) ? 4044 : (x < 16**14) ? 4040 : (x < 16**15) ? 4036 : (x < 16**16) ? 4032 : (x < 16**17) ? 4028 : (x < 16**18) ? 4024 : (x < 16**19) ? 4020 : (x < 16**20) ? 4016 : (x < 16**21) ? 4012 : (x < 16**22) ? 4008 : (x < 16**23) ? 4004 : (x < 16**24) ? 4000 : (x < 16**25) ? 3996 : (x < 16**26) ? 3992 : (x < 16**27) ? 3988 : (x < 16**28) ? 3984 : (x < 16**29) ? 3980 : (x < 16**30) ? 3976 : (x < 16**31) ? 3972 : (x < 16**32) ? 3968 : (x < 16**33) ? 3964 : (x < 16**34) ? 3960 : (x < 16**35) ? 3956 : (x < 16**36) ? 3952 : (x < 16**37) ? 3948 : (x < 16**38) ? 3944 : (x < 16**39) ? 3940 : (x < 16**40) ? 3936 : (x < 16**41) ? 3932 : (x < 16**42) ? 3928 : (x < 16**43) ? 3924 : (x < 16**44) ? 3920 : (x < 16**45) ? 3916 : (x < 16**46) ? 3912 : (x < 16**47) ? 3908 : (x < 16**48) ? 3904 : (x < 16**49) ? 3900 : (x < 16**50) ? 3896 : (x < 16**51) ? 3892 : (x < 16**52) ? 3888 : (x < 16**53) ? 3884 : (x < 16**54) ? 3880 : (x < 16**55) ? 3876 : (x < 16**56) ? 3872 : (x < 16**57) ? 3868 : (x < 16**58) ? 3864 : (x < 16**59) ? 3860 : (x < 16**60) ? 3856 : (x < 16**61) ? 3852 : (x < 16**62) ? 3848 : (x < 16**63) ? 3844 : (x < 16**64) ? 3840 : (x < 16**65) ? 3836 : (x < 16**66) ? 3832 : (x < 16**67) ? 3828 : (x < 16**68) ? 3824 : (x < 16**69) ? 3820 : (x < 16**70) ? 3816 : (x < 16**71) ? 3812 : (x < 16**72) ? 3808 : (x < 16**73) ? 3804 : (x < 16**74) ? 3800 : (x < 16**75) ? 3796 : (x < 16**76) ? 3792 : (x < 16**77) ? 3788 : (x < 16**78) ? 3784 : (x < 16**79) ? 3780 : (x < 16**80) ? 3776 : (x < 16**81) ? 3772 : (x < 16**82) ? 3768 : (x < 16**83) ? 3764 : (x < 16**84) ? 3760 : (x < 16**85) ? 3756 : (x < 16**86) ? 3752 : (x < 16**87) ? 3748 : (x < 16**88) ? 3744 : (x < 16**89) ? 3740 : (x < 16**90) ? 3736 : (x < 16**91) ? 3732 : (x < 16**92) ? 3728 : (x < 16**93) ? 3724 : (x < 16**94) ? 3720 : (x < 16**95) ? 3716 : (x < 16**96) ? 3712 : (x < 16**97) ? 3708 : (x < 16**98) ? 3704 : (x < 16**99) ? 3700 : (x < 16**100) ? 3696 : (x < 16**101) ? 3692 : (x < 16**102) ? 3688 : (x < 16**103) ? 3684 : (x < 16**104) ? 3680 : (x < 16**105) ? 3676 : (x < 16**106) ? 3672 : (x < 16**107) ? 3668 : (x < 16**108) ? 3664 : (x < 16**109) ? 3660 : (x < 16**110) ? 3656 : (x < 16**111) ? 3652 : (x < 16**112) ? 3648 : (x < 16**113) ? 3644 : (x < 16**114) ? 3640 : (x < 16**115) ? 3636 : (x < 16**116) ? 3632 : (x < 16**117) ? 3628 : (x < 16**118) ? 3624 : (x < 16**119) ? 3620 : (x < 16**120) ? 3616 : (x < 16**121) ? 3612 : (x < 16**122) ? 3608 : (x < 16**123) ? 3604 : (x < 16**124) ? 3600 : (x < 16**125) ? 3596 : (x < 16**126) ? 3592 : (x < 16**127) ? 3588 : (x < 16**128) ? 3584 : (x < 16**129) ? 3580 : (x < 16**130) ? 3576 : (x < 16**131) ? 3572 : (x < 16**132) ? 3568 : (x < 16**133) ? 3564 : (x < 16**134) ? 3560 : (x < 16**135) ? 3556 : (x < 16**136) ? 3552 : (x < 16**137) ? 3548 : (x < 16**138) ? 3544 : (x < 16**139) ? 3540 : (x < 16**140) ? 3536 : (x < 16**141) ? 3532 : (x < 16**142) ? 3528 : (x < 16**143) ? 3524 : (x < 16**144) ? 3520 : (x < 16**145) ? 3516 : (x < 16**146) ? 3512 : (x < 16**147) ? 3508 : (x < 16**148) ? 3504 : (x < 16**149) ? 3500 : (x < 16**150) ? 3496 : (x < 16**151) ? 3492 : (x < 16**152) ? 3488 : (x < 16**153) ? 3484 : (x < 16**154) ? 3480 : (x < 16**155) ? 3476 : (x < 16**156) ? 3472 : (x < 16**157) ? 3468 : (x < 16**158) ? 3464 : (x < 16**159) ? 3460 : (x < 16**160) ? 3456 : (x < 16**161) ? 3452 : (x < 16**162) ? 3448 : (x < 16**163) ? 3444 : (x < 16**164) ? 3440 : (x < 16**165) ? 3436 : (x < 16**166) ? 3432 : (x < 16**167) ? 3428 : (x < 16**168) ? 3424 : (x < 16**169) ? 3420 : (x < 16**170) ? 3416 : (x < 16**171) ? 3412 : (x < 16**172) ? 3408 : (x < 16**173) ? 3404 : (x < 16**174) ? 3400 : (x < 16**175) ? 3396 : (x < 16**176) ? 3392 : (x < 16**177) ? 3388 : (x < 16**178) ? 3384 : (x < 16**179) ? 3380 : (x < 16**180) ? 3376 : (x < 16**181) ? 3372 : (x < 16**182) ? 3368 : (x < 16**183) ? 3364 : (x < 16**184) ? 3360 : (x < 16**185) ? 3356 : (x < 16**186) ? 3352 : (x < 16**187) ? 3348 : (x < 16**188) ? 3344 : (x < 16**189) ? 3340 : (x < 16**190) ? 3336 : (x < 16**191) ? 3332 : (x < 16**192) ? 3328 : (x < 16**193) ? 3324 : (x < 16**194) ? 3320 : (x < 16**195) ? 3316 : (x < 16**196) ? 3312 : (x < 16**197) ? 3308 : (x < 16**198) ? 3304 : (x < 16**199) ? 3300 : (x < 16**200) ? 3296 : (x < 16**201) ? 3292 : (x < 16**202) ? 3288 : (x < 16**203) ? 3284 : (x < 16**204) ? 3280 : (x < 16**205) ? 3276 : (x < 16**206) ? 3272 : (x < 16**207) ? 3268 : (x < 16**208) ? 3264 : (x < 16**209) ? 3260 : (x < 16**210) ? 3256 : (x < 16**211) ? 3252 : (x < 16**212) ? 3248 : (x < 16**213) ? 3244 : (x < 16**214) ? 3240 : (x < 16**215) ? 3236 : (x < 16**216) ? 3232 : (x < 16**217) ? 3228 : (x < 16**218) ? 3224 : (x < 16**219) ? 3220 : (x < 16**220) ? 3216 : (x < 16**221) ? 3212 : (x < 16**222) ? 3208 : (x < 16**223) ? 3204 : (x < 16**224) ? 3200 : (x < 16**225) ? 3196 : (x < 16**226) ? 3192 : (x < 16**227) ? 3188 : (x < 16**228) ? 3184 : (x < 16**229) ? 3180 : (x < 16**230) ? 3176 : (x < 16**231) ? 3172 : (x < 16**232) ? 3168 : (x < 16**233) ? 3164 : (x < 16**234) ? 3160 : (x < 16**235) ? 3156 : (x < 16**236) ? 3152 : (x < 16**237) ? 3148 : (x < 16**238) ? 3144 : (x < 16**239) ? 3140 : (x < 16**240) ? 3136 : (x < 16**241) ? 3132 : (x < 16**242) ? 3128 : (x < 16**243) ? 3124 : (x < 16**244) ? 3120 : (x < 16**245) ? 3116 : (x < 16**246) ? 3112 : (x < 16**247) ? 3108 : (x < 16**248) ? 3104 : (x < 16**249) ? 3100 : (x < 16**250) ? 3096 : (x < 16**251) ? 3092 : (x < 16**252) ? 3088 : (x < 16**253) ? 3084 : (x < 16**254) ? 3080 : (x < 16**255) ? 3076 : (x < 16**256) ? 3072 : (x < 16**257) ? 3068 : (x < 16**258) ? 3064 : (x < 16**259) ? 3060 : (x < 16**260) ? 3056 : (x < 16**261) ? 3052 : (x < 16**262) ? 3048 : (x < 16**263) ? 3044 : (x < 16**264) ? 3040 : (x < 16**265) ? 3036 : (x < 16**266) ? 3032 : (x < 16**267) ? 3028 : (x < 16**268) ? 3024 : (x < 16**269) ? 3020 : (x < 16**270) ? 3016 : (x < 16**271) ? 3012 : (x < 16**272) ? 3008 : (x < 16**273) ? 3004 : (x < 16**274) ? 3000 : (x < 16**275) ? 2996 : (x < 16**276) ? 2992 : (x < 16**277) ? 2988 : (x < 16**278) ? 2984 : (x < 16**279) ? 2980 : (x < 16**280) ? 2976 : (x < 16**281) ? 2972 : (x < 16**282) ? 2968 : (x < 16**283) ? 2964 : (x < 16**284) ? 2960 : (x < 16**285) ? 2956 : (x < 16**286) ? 2952 : (x < 16**287) ? 2948 : (x < 16**288) ? 2944 : (x < 16**289) ? 2940 : (x < 16**290) ? 2936 : (x < 16**291) ? 2932 : (x < 16**292) ? 2928 : (x < 16**293) ? 2924 : (x < 16**294) ? 2920 : (x < 16**295) ? 2916 : (x < 16**296) ? 2912 : (x < 16**297) ? 2908 : (x < 16**298) ? 2904 : (x < 16**299) ? 2900 : (x < 16**300) ? 2896 : (x < 16**301) ? 2892 : (x < 16**302) ? 2888 : (x < 16**303) ? 2884 : (x < 16**304) ? 2880 : (x < 16**305) ? 2876 : (x < 16**306) ? 2872 : (x < 16**307) ? 2868 : (x < 16**308) ? 2864 : (x < 16**309) ? 2860 : (x < 16**310) ? 2856 : (x < 16**311) ? 2852 : (x < 16**312) ? 2848 : (x < 16**313) ? 2844 : (x < 16**314) ? 2840 : (x < 16**315) ? 2836 : (x < 16**316) ? 2832 : (x < 16**317) ? 2828 : (x < 16**318) ? 2824 : (x < 16**319) ? 2820 : (x < 16**320) ? 2816 : (x < 16**321) ? 2812 : (x < 16**322) ? 2808 : (x < 16**323) ? 2804 : (x < 16**324) ? 2800 : (x < 16**325) ? 2796 : (x < 16**326) ? 2792 : (x < 16**327) ? 2788 : (x < 16**328) ? 2784 : (x < 16**329) ? 2780 : (x < 16**330) ? 2776 : (x < 16**331) ? 2772 : (x < 16**332) ? 2768 : (x < 16**333) ? 2764 : (x < 16**334) ? 2760 : (x < 16**335) ? 2756 : (x < 16**336) ? 2752 : (x < 16**337) ? 2748 : (x < 16**338) ? 2744 : (x < 16**339) ? 2740 : (x < 16**340) ? 2736 : (x < 16**341) ? 2732 : (x < 16**342) ? 2728 : (x < 16**343) ? 2724 : (x < 16**344) ? 2720 : (x < 16**345) ? 2716 : (x < 16**346) ? 2712 : (x < 16**347) ? 2708 : (x < 16**348) ? 2704 : (x < 16**349) ? 2700 : (x < 16**350) ? 2696 : (x < 16**351) ? 2692 : (x < 16**352) ? 2688 : (x < 16**353) ? 2684 : (x < 16**354) ? 2680 : (x < 16**355) ? 2676 : (x < 16**356) ? 2672 : (x < 16**357) ? 2668 : (x < 16**358) ? 2664 : (x < 16**359) ? 2660 : (x < 16**360) ? 2656 : (x < 16**361) ? 2652 : (x < 16**362) ? 2648 : (x < 16**363) ? 2644 : (x < 16**364) ? 2640 : (x < 16**365) ? 2636 : (x < 16**366) ? 2632 : (x < 16**367) ? 2628 : (x < 16**368) ? 2624 : (x < 16**369) ? 2620 : (x < 16**370) ? 2616 : (x < 16**371) ? 2612 : (x < 16**372) ? 2608 : (x < 16**373) ? 2604 : (x < 16**374) ? 2600 : (x < 16**375) ? 2596 : (x < 16**376) ? 2592 : (x < 16**377) ? 2588 : (x < 16**378) ? 2584 : (x < 16**379) ? 2580 : (x < 16**380) ? 2576 : (x < 16**381) ? 2572 : (x < 16**382) ? 2568 : (x < 16**383) ? 2564 : (x < 16**384) ? 2560 : (x < 16**385) ? 2556 : (x < 16**386) ? 2552 : (x < 16**387) ? 2548 : (x < 16**388) ? 2544 : (x < 16**389) ? 2540 : (x < 16**390) ? 2536 : (x < 16**391) ? 2532 : (x < 16**392) ? 2528 : (x < 16**393) ? 2524 : (x < 16**394) ? 2520 : (x < 16**395) ? 2516 : (x < 16**396) ? 2512 : (x < 16**397) ? 2508 : (x < 16**398) ? 2504 : (x < 16**399) ? 2500 : (x < 16**400) ? 2496 : (x < 16**401) ? 2492 : (x < 16**402) ? 2488 : (x < 16**403) ? 2484 : (x < 16**404) ? 2480 : (x < 16**405) ? 2476 : (x < 16**406) ? 2472 : (x < 16**407) ? 2468 : (x < 16**408) ? 2464 : (x < 16**409) ? 2460 : (x < 16**410) ? 2456 : (x < 16**411) ? 2452 : (x < 16**412) ? 2448 : (x < 16**413) ? 2444 : (x < 16**414) ? 2440 : (x < 16**415) ? 2436 : (x < 16**416) ? 2432 : (x < 16**417) ? 2428 : (x < 16**418) ? 2424 : (x < 16**419) ? 2420 : (x < 16**420) ? 2416 : (x < 16**421) ? 2412 : (x < 16**422) ? 2408 : (x < 16**423) ? 2404 : (x < 16**424) ? 2400 : (x < 16**425) ? 2396 : (x < 16**426) ? 2392 : (x < 16**427) ? 2388 : (x < 16**428) ? 2384 : (x < 16**429) ? 2380 : (x < 16**430) ? 2376 : (x < 16**431) ? 2372 : (x < 16**432) ? 2368 : (x < 16**433) ? 2364 : (x < 16**434) ? 2360 : (x < 16**435) ? 2356 : (x < 16**436) ? 2352 : (x < 16**437) ? 2348 : (x < 16**438) ? 2344 : (x < 16**439) ? 2340 : (x < 16**440) ? 2336 : (x < 16**441) ? 2332 : (x < 16**442) ? 2328 : (x < 16**443) ? 2324 : (x < 16**444) ? 2320 : (x < 16**445) ? 2316 : (x < 16**446) ? 2312 : (x < 16**447) ? 2308 : (x < 16**448) ? 2304 : (x < 16**449) ? 2300 : (x < 16**450) ? 2296 : (x < 16**451) ? 2292 : (x < 16**452) ? 2288 : (x < 16**453) ? 2284 : (x < 16**454) ? 2280 : (x < 16**455) ? 2276 : (x < 16**456) ? 2272 : (x < 16**457) ? 2268 : (x < 16**458) ? 2264 : (x < 16**459) ? 2260 : (x < 16**460) ? 2256 : (x < 16**461) ? 2252 : (x < 16**462) ? 2248 : (x < 16**463) ? 2244 : (x < 16**464) ? 2240 : (x < 16**465) ? 2236 : (x < 16**466) ? 2232 : (x < 16**467) ? 2228 : (x < 16**468) ? 2224 : (x < 16**469) ? 2220 : (x < 16**470) ? 2216 : (x < 16**471) ? 2212 : (x < 16**472) ? 2208 : (x < 16**473) ? 2204 : (x < 16**474) ? 2200 : (x < 16**475) ? 2196 : (x < 16**476) ? 2192 : (x < 16**477) ? 2188 : (x < 16**478) ? 2184 : (x < 16**479) ? 2180 : (x < 16**480) ? 2176 : (x < 16**481) ? 2172 : (x < 16**482) ? 2168 : (x < 16**483) ? 2164 : (x < 16**484) ? 2160 : (x < 16**485) ? 2156 : (x < 16**486) ? 2152 : (x < 16**487) ? 2148 : (x < 16**488) ? 2144 : (x < 16**489) ? 2140 : (x < 16**490) ? 2136 : (x < 16**491) ? 2132 : (x < 16**492) ? 2128 : (x < 16**493) ? 2124 : (x < 16**494) ? 2120 : (x < 16**495) ? 2116 : (x < 16**496) ? 2112 : (x < 16**497) ? 2108 : (x < 16**498) ? 2104 : (x < 16**499) ? 2100 : (x < 16**500) ? 2096 : (x < 16**501) ? 2092 : (x < 16**502) ? 2088 : (x < 16**503) ? 2084 : (x < 16**504) ? 2080 : (x < 16**505) ? 2076 : (x < 16**506) ? 2072 : (x < 16**507) ? 2068 : (x < 16**508) ? 2064 : (x < 16**509) ? 2060 : (x < 16**510) ? 2056 : (x < 16**511) ? 2052 : (x < 16**512) ? 2048 : (x < 16**513) ? 2044 : (x < 16**514) ? 2040 : (x < 16**515) ? 2036 : (x < 16**516) ? 2032 : (x < 16**517) ? 2028 : (x < 16**518) ? 2024 : (x < 16**519) ? 2020 : (x < 16**520) ? 2016 : (x < 16**521) ? 2012 : (x < 16**522) ? 2008 : (x < 16**523) ? 2004 : (x < 16**524) ? 2000 : (x < 16**525) ? 1996 : (x < 16**526) ? 1992 : (x < 16**527) ? 1988 : (x < 16**528) ? 1984 : (x < 16**529) ? 1980 : (x < 16**530) ? 1976 : (x < 16**531) ? 1972 : (x < 16**532) ? 1968 : (x < 16**533) ? 1964 : (x < 16**534) ? 1960 : (x < 16**535) ? 1956 : (x < 16**536) ? 1952 : (x < 16**537) ? 1948 : (x < 16**538) ? 1944 : (x < 16**539) ? 1940 : (x < 16**540) ? 1936 : (x < 16**541) ? 1932 : (x < 16**542) ? 1928 : (x < 16**543) ? 1924 : (x < 16**544) ? 1920 : (x < 16**545) ? 1916 : (x < 16**546) ? 1912 : (x < 16**547) ? 1908 : (x < 16**548) ? 1904 : (x < 16**549) ? 1900 : (x < 16**550) ? 1896 : (x < 16**551) ? 1892 : (x < 16**552) ? 1888 : (x < 16**553) ? 1884 : (x < 16**554) ? 1880 : (x < 16**555) ? 1876 : (x < 16**556) ? 1872 : (x < 16**557) ? 1868 : (x < 16**558) ? 1864 : (x < 16**559) ? 1860 : (x < 16**560) ? 1856 : (x < 16**561) ? 1852 : (x < 16**562) ? 1848 : (x < 16**563) ? 1844 : (x < 16**564) ? 1840 : (x < 16**565) ? 1836 : (x < 16**566) ? 1832 : (x < 16**567) ? 1828 : (x < 16**568) ? 1824 : (x < 16**569) ? 1820 : (x < 16**570) ? 1816 : (x < 16**571) ? 1812 : (x < 16**572) ? 1808 : (x < 16**573) ? 1804 : (x < 16**574) ? 1800 : (x < 16**575) ? 1796 : (x < 16**576) ? 1792 : (x < 16**577) ? 1788 : (x < 16**578) ? 1784 : (x < 16**579) ? 1780 : (x < 16**580) ? 1776 : (x < 16**581) ? 1772 : (x < 16**582) ? 1768 : (x < 16**583) ? 1764 : (x < 16**584) ? 1760 : (x < 16**585) ? 1756 : (x < 16**586) ? 1752 : (x < 16**587) ? 1748 : (x < 16**588) ? 1744 : (x < 16**589) ? 1740 : (x < 16**590) ? 1736 : (x < 16**591) ? 1732 : (x < 16**592) ? 1728 : (x < 16**593) ? 1724 : (x < 16**594) ? 1720 : (x < 16**595) ? 1716 : (x < 16**596) ? 1712 : (x < 16**597) ? 1708 : (x < 16**598) ? 1704 : (x < 16**599) ? 1700 : (x < 16**600) ? 1696 : (x < 16**601) ? 1692 : (x < 16**602) ? 1688 : (x < 16**603) ? 1684 : (x < 16**604) ? 1680 : (x < 16**605) ? 1676 : (x < 16**606) ? 1672 : (x < 16**607) ? 1668 : (x < 16**608) ? 1664 : (x < 16**609) ? 1660 : (x < 16**610) ? 1656 : (x < 16**611) ? 1652 : (x < 16**612) ? 1648 : (x < 16**613) ? 1644 : (x < 16**614) ? 1640 : (x < 16**615) ? 1636 : (x < 16**616) ? 1632 : (x < 16**617) ? 1628 : (x < 16**618) ? 1624 : (x < 16**619) ? 1620 : (x < 16**620) ? 1616 : (x < 16**621) ? 1612 : (x < 16**622) ? 1608 : (x < 16**623) ? 1604 : (x < 16**624) ? 1600 : (x < 16**625) ? 1596 : (x < 16**626) ? 1592 : (x < 16**627) ? 1588 : (x < 16**628) ? 1584 : (x < 16**629) ? 1580 : (x < 16**630) ? 1576 : (x < 16**631) ? 1572 : (x < 16**632) ? 1568 : (x < 16**633) ? 1564 : (x < 16**634) ? 1560 : (x < 16**635) ? 1556 : (x < 16**636) ? 1552 : (x < 16**637) ? 1548 : (x < 16**638) ? 1544 : (x < 16**639) ? 1540 : (x < 16**640) ? 1536 : (x < 16**641) ? 1532 : (x < 16**642) ? 1528 : (x < 16**643) ? 1524 : (x < 16**644) ? 1520 : (x < 16**645) ? 1516 : (x < 16**646) ? 1512 : (x < 16**647) ? 1508 : (x < 16**648) ? 1504 : (x < 16**649) ? 1500 : (x < 16**650) ? 1496 : (x < 16**651) ? 1492 : (x < 16**652) ? 1488 : (x < 16**653) ? 1484 : (x < 16**654) ? 1480 : (x < 16**655) ? 1476 : (x < 16**656) ? 1472 : (x < 16**657) ? 1468 : (x < 16**658) ? 1464 : (x < 16**659) ? 1460 : (x < 16**660) ? 1456 : (x < 16**661) ? 1452 : (x < 16**662) ? 1448 : (x < 16**663) ? 1444 : (x < 16**664) ? 1440 : (x < 16**665) ? 1436 : (x < 16**666) ? 1432 : (x < 16**667) ? 1428 : (x < 16**668) ? 1424 : (x < 16**669) ? 1420 : (x < 16**670) ? 1416 : (x < 16**671) ? 1412 : (x < 16**672) ? 1408 : (x < 16**673) ? 1404 : (x < 16**674) ? 1400 : (x < 16**675) ? 1396 : (x < 16**676) ? 1392 : (x < 16**677) ? 1388 : (x < 16**678) ? 1384 : (x < 16**679) ? 1380 : (x < 16**680) ? 1376 : (x < 16**681) ? 1372 : (x < 16**682) ? 1368 : (x < 16**683) ? 1364 : (x < 16**684) ? 1360 : (x < 16**685) ? 1356 : (x < 16**686) ? 1352 : (x < 16**687) ? 1348 : (x < 16**688) ? 1344 : (x < 16**689) ? 1340 : (x < 16**690) ? 1336 : (x < 16**691) ? 1332 : (x < 16**692) ? 1328 : (x < 16**693) ? 1324 : (x < 16**694) ? 1320 : (x < 16**695) ? 1316 : (x < 16**696) ? 1312 : (x < 16**697) ? 1308 : (x < 16**698) ? 1304 : (x < 16**699) ? 1300 : (x < 16**700) ? 1296 : (x < 16**701) ? 1292 : (x < 16**702) ? 1288 : (x < 16**703) ? 1284 : (x < 16**704) ? 1280 : (x < 16**705) ? 1276 : (x < 16**706) ? 1272 : (x < 16**707) ? 1268 : (x < 16**708) ? 1264 : (x < 16**709) ? 1260 : (x < 16**710) ? 1256 : (x < 16**711) ? 1252 : (x < 16**712) ? 1248 : (x < 16**713) ? 1244 : (x < 16**714) ? 1240 : (x < 16**715) ? 1236 : (x < 16**716) ? 1232 : (x < 16**717) ? 1228 : (x < 16**718) ? 1224 : (x < 16**719) ? 1220 : (x < 16**720) ? 1216 : (x < 16**721) ? 1212 : (x < 16**722) ? 1208 : (x < 16**723) ? 1204 : (x < 16**724) ? 1200 : (x < 16**725) ? 1196 : (x < 16**726) ? 1192 : (x < 16**727) ? 1188 : (x < 16**728) ? 1184 : (x < 16**729) ? 1180 : (x < 16**730) ? 1176 : (x < 16**731) ? 1172 : (x < 16**732) ? 1168 : (x < 16**733) ? 1164 : (x < 16**734) ? 1160 : (x < 16**735) ? 1156 : (x < 16**736) ? 1152 : (x < 16**737) ? 1148 : (x < 16**738) ? 1144 : (x < 16**739) ? 1140 : (x < 16**740) ? 1136 : (x < 16**741) ? 1132 : (x < 16**742) ? 1128 : (x < 16**743) ? 1124 : (x < 16**744) ? 1120 : (x < 16**745) ? 1116 : (x < 16**746) ? 1112 : (x < 16**747) ? 1108 : (x < 16**748) ? 1104 : (x < 16**749) ? 1100 : (x < 16**750) ? 1096 : (x < 16**751) ? 1092 : (x < 16**752) ? 1088 : (x < 16**753) ? 1084 : (x < 16**754) ? 1080 : (x < 16**755) ? 1076 : (x < 16**756) ? 1072 : (x < 16**757) ? 1068 : (x < 16**758) ? 1064 : (x < 16**759) ? 1060 : (x < 16**760) ? 1056 : (x < 16**761) ? 1052 : (x < 16**762) ? 1048 : (x < 16**763) ? 1044 : (x < 16**764) ? 1040 : (x < 16**765) ? 1036 : (x < 16**766) ? 1032 : (x < 16**767) ? 1028 : (x < 16**768) ? 1024 : (x < 16**769) ? 1020 : (x < 16**770) ? 1016 : (x < 16**771) ? 1012 : (x < 16**772) ? 1008 : (x < 16**773) ? 1004 : (x < 16**774) ? 1000 : (x < 16**775) ? 996 : (x < 16**776) ? 992 : (x < 16**777) ? 988 : (x < 16**778) ? 984 : (x < 16**779) ? 980 : (x < 16**780) ? 976 : (x < 16**781) ? 972 : (x < 16**782) ? 968 : (x < 16**783) ? 964 : (x < 16**784) ? 960 : (x < 16**785) ? 956 : (x < 16**786) ? 952 : (x < 16**787) ? 948 : (x < 16**788) ? 944 : (x < 16**789) ? 940 : (x < 16**790) ? 936 : (x < 16**791) ? 932 : (x < 16**792) ? 928 : (x < 16**793) ? 924 : (x < 16**794) ? 920 : (x < 16**795) ? 916 : (x < 16**796) ? 912 : (x < 16**797) ? 908 : (x < 16**798) ? 904 : (x < 16**799) ? 900 : (x < 16**800) ? 896 : (x < 16**801) ? 892 : (x < 16**802) ? 888 : (x < 16**803) ? 884 : (x < 16**804) ? 880 : (x < 16**805) ? 876 : (x < 16**806) ? 872 : (x < 16**807) ? 868 : (x < 16**808) ? 864 : (x < 16**809) ? 860 : (x < 16**810) ? 856 : (x < 16**811) ? 852 : (x < 16**812) ? 848 : (x < 16**813) ? 844 : (x < 16**814) ? 840 : (x < 16**815) ? 836 : (x < 16**816) ? 832 : (x < 16**817) ? 828 : (x < 16**818) ? 824 : (x < 16**819) ? 820 : (x < 16**820) ? 816 : (x < 16**821) ? 812 : (x < 16**822) ? 808 : (x < 16**823) ? 804 : (x < 16**824) ? 800 : (x < 16**825) ? 796 : (x < 16**826) ? 792 : (x < 16**827) ? 788 : (x < 16**828) ? 784 : (x < 16**829) ? 780 : (x < 16**830) ? 776 : (x < 16**831) ? 772 : (x < 16**832) ? 768 : (x < 16**833) ? 764 : (x < 16**834) ? 760 : (x < 16**835) ? 756 : (x < 16**836) ? 752 : (x < 16**837) ? 748 : (x < 16**838) ? 744 : (x < 16**839) ? 740 : (x < 16**840) ? 736 : (x < 16**841) ? 732 : (x < 16**842) ? 728 : (x < 16**843) ? 724 : (x < 16**844) ? 720 : (x < 16**845) ? 716 : (x < 16**846) ? 712 : (x < 16**847) ? 708 : (x < 16**848) ? 704 : (x < 16**849) ? 700 : (x < 16**850) ? 696 : (x < 16**851) ? 692 : (x < 16**852) ? 688 : (x < 16**853) ? 684 : (x < 16**854) ? 680 : (x < 16**855) ? 676 : (x < 16**856) ? 672 : (x < 16**857) ? 668 : (x < 16**858) ? 664 : (x < 16**859) ? 660 : (x < 16**860) ? 656 : (x < 16**861) ? 652 : (x < 16**862) ? 648 : (x < 16**863) ? 644 : (x < 16**864) ? 640 : (x < 16**865) ? 636 : (x < 16**866) ? 632 : (x < 16**867) ? 628 : (x < 16**868) ? 624 : (x < 16**869) ? 620 : (x < 16**870) ? 616 : (x < 16**871) ? 612 : (x < 16**872) ? 608 : (x < 16**873) ? 604 : (x < 16**874) ? 600 : (x < 16**875) ? 596 : (x < 16**876) ? 592 : (x < 16**877) ? 588 : (x < 16**878) ? 584 : (x < 16**879) ? 580 : (x < 16**880) ? 576 : (x < 16**881) ? 572 : (x < 16**882) ? 568 : (x < 16**883) ? 564 : (x < 16**884) ? 560 : (x < 16**885) ? 556 : (x < 16**886) ? 552 : (x < 16**887) ? 548 : (x < 16**888) ? 544 : (x < 16**889) ? 540 : (x < 16**890) ? 536 : (x < 16**891) ? 532 : (x < 16**892) ? 528 : (x < 16**893) ? 524 : (x < 16**894) ? 520 : (x < 16**895) ? 516 : (x < 16**896) ? 512 : (x < 16**897) ? 508 : (x < 16**898) ? 504 : (x < 16**899) ? 500 : (x < 16**900) ? 496 : (x < 16**901) ? 492 : (x < 16**902) ? 488 : (x < 16**903) ? 484 : (x < 16**904) ? 480 : (x < 16**905) ? 476 : (x < 16**906) ? 472 : (x < 16**907) ? 468 : (x < 16**908) ? 464 : (x < 16**909) ? 460 : (x < 16**910) ? 456 : (x < 16**911) ? 452 : (x < 16**912) ? 448 : (x < 16**913) ? 444 : (x < 16**914) ? 440 : (x < 16**915) ? 436 : (x < 16**916) ? 432 : (x < 16**917) ? 428 : (x < 16**918) ? 424 : (x < 16**919) ? 420 : (x < 16**920) ? 416 : (x < 16**921) ? 412 : (x < 16**922) ? 408 : (x < 16**923) ? 404 : (x < 16**924) ? 400 : (x < 16**925) ? 396 : (x < 16**926) ? 392 : (x < 16**927) ? 388 : (x < 16**928) ? 384 : (x < 16**929) ? 380 : (x < 16**930) ? 376 : (x < 16**931) ? 372 : (x < 16**932) ? 368 : (x < 16**933) ? 364 : (x < 16**934) ? 360 : (x < 16**935) ? 356 : (x < 16**936) ? 352 : (x < 16**937) ? 348 : (x < 16**938) ? 344 : (x < 16**939) ? 340 : (x < 16**940) ? 336 : (x < 16**941) ? 332 : (x < 16**942) ? 328 : (x < 16**943) ? 324 : (x < 16**944) ? 320 : (x < 16**945) ? 316 : (x < 16**946) ? 312 : (x < 16**947) ? 308 : (x < 16**948) ? 304 : (x < 16**949) ? 300 : (x < 16**950) ? 296 : (x < 16**951) ? 292 : (x < 16**952) ? 288 : (x < 16**953) ? 284 : (x < 16**954) ? 280 : (x < 16**955) ? 276 : (x < 16**956) ? 272 : (x < 16**957) ? 268 : (x < 16**958) ? 264 : (x < 16**959) ? 260 : (x < 16**960) ? 256 : (x < 16**961) ? 252 : (x < 16**962) ? 248 : (x < 16**963) ? 244 : (x < 16**964) ? 240 : (x < 16**965) ? 236 : (x < 16**966) ? 232 : (x < 16**967) ? 228 : (x < 16**968) ? 224 : (x < 16**969) ? 220 : (x < 16**970) ? 216 : (x < 16**971) ? 212 : (x < 16**972) ? 208 : (x < 16**973) ? 204 : (x < 16**974) ? 200 : (x < 16**975) ? 196 : (x < 16**976) ? 192 : (x < 16**977) ? 188 : (x < 16**978) ? 184 : (x < 16**979) ? 180 : (x < 16**980) ? 176 : (x < 16**981) ? 172 : (x < 16**982) ? 168 : (x < 16**983) ? 164 : (x < 16**984) ? 160 : (x < 16**985) ? 156 : (x < 16**986) ? 152 : (x < 16**987) ? 148 : (x < 16**988) ? 144 : (x < 16**989) ? 140 : (x < 16**990) ? 136 : (x < 16**991) ? 132 : (x < 16**992) ? 128 : (x < 16**993) ? 124 : (x < 16**994) ? 120 : (x < 16**995) ? 116 : (x < 16**996) ? 112 : (x < 16**997) ? 108 : (x < 16**998) ? 104 : (x < 16**999) ? 100 : (x < 16**1000) ? 96 : (x < 16**1001) ? 92 : (x < 16**1002) ? 88 : (x < 16**1003) ? 84 : (x < 16**1004) ? 80 : (x < 16**1005) ? 76 : (x < 16**1006) ? 72 : (x < 16**1007) ? 68 : (x < 16**1008) ? 64 : (x < 16**1009) ? 60 : (x < 16**1010) ? 56 : (x < 16**1011) ? 52 : (x < 16**1012) ? 48 : (x < 16**1013) ? 44 : (x < 16**1014) ? 40 : (x < 16**1015) ? 36 : (x < 16**1016) ? 32 : (x < 16**1017) ? 28 : (x < 16**1018) ? 24 : (x < 16**1019) ? 20 : (x < 16**1020) ? 16 : (x < 16**1021) ? 12 : (x < 16**1022) ? 8 : (x < 16**1023) ? 4 : (x < 16**1024) ? 0 : 0


`define rotate(x)\
{x[4039:4032],x[4047:4040],x[4055:4048],x[4063:4056],x[4071:4064],x[4079:4072],x[4087:4080],x[4095:4088],x[3975:3968],x[3983:3976],x[3991:3984],x[3999:3992],x[4007:4000],x[4015:4008],x[4023:4016],x[4031:4024],x[3911:3904],x[3919:3912],x[3927:3920],x[3935:3928],x[3943:3936],x[3951:3944],x[3959:3952],x[3967:3960],x[3847:3840],x[3855:3848],x[3863:3856],x[3871:3864],x[3879:3872],x[3887:3880],x[3895:3888],x[3903:3896],x[3783:3776],x[3791:3784],x[3799:3792],x[3807:3800],x[3815:3808],x[3823:3816],x[3831:3824],x[3839:3832],x[3719:3712],x[3727:3720],x[3735:3728],x[3743:3736],x[3751:3744],x[3759:3752],x[3767:3760],x[3775:3768],x[3655:3648],x[3663:3656],x[3671:3664],x[3679:3672],x[3687:3680],x[3695:3688],x[3703:3696],x[3711:3704],x[3591:3584],x[3599:3592],x[3607:3600],x[3615:3608],x[3623:3616],x[3631:3624],x[3639:3632],x[3647:3640],x[3527:3520],x[3535:3528],x[3543:3536],x[3551:3544],x[3559:3552],x[3567:3560],x[3575:3568],x[3583:3576],x[3463:3456],x[3471:3464],x[3479:3472],x[3487:3480],x[3495:3488],x[3503:3496],x[3511:3504],x[3519:3512],x[3399:3392],x[3407:3400],x[3415:3408],x[3423:3416],x[3431:3424],x[3439:3432],x[3447:3440],x[3455:3448],x[3335:3328],x[3343:3336],x[3351:3344],x[3359:3352],x[3367:3360],x[3375:3368],x[3383:3376],x[3391:3384],x[3271:3264],x[3279:3272],x[3287:3280],x[3295:3288],x[3303:3296],x[3311:3304],x[3319:3312],x[3327:3320],x[3207:3200],x[3215:3208],x[3223:3216],x[3231:3224],x[3239:3232],x[3247:3240],x[3255:3248],x[3263:3256],x[3143:3136],x[3151:3144],x[3159:3152],x[3167:3160],x[3175:3168],x[3183:3176],x[3191:3184],x[3199:3192],x[3079:3072],x[3087:3080],x[3095:3088],x[3103:3096],x[3111:3104],x[3119:3112],x[3127:3120],x[3135:3128],x[3015:3008],x[3023:3016],x[3031:3024],x[3039:3032],x[3047:3040],x[3055:3048],x[3063:3056],x[3071:3064],x[2951:2944],x[2959:2952],x[2967:2960],x[2975:2968],x[2983:2976],x[2991:2984],x[2999:2992],x[3007:3000],x[2887:2880],x[2895:2888],x[2903:2896],x[2911:2904],x[2919:2912],x[2927:2920],x[2935:2928],x[2943:2936],x[2823:2816],x[2831:2824],x[2839:2832],x[2847:2840],x[2855:2848],x[2863:2856],x[2871:2864],x[2879:2872],x[2759:2752],x[2767:2760],x[2775:2768],x[2783:2776],x[2791:2784],x[2799:2792],x[2807:2800],x[2815:2808],x[2695:2688],x[2703:2696],x[2711:2704],x[2719:2712],x[2727:2720],x[2735:2728],x[2743:2736],x[2751:2744],x[2631:2624],x[2639:2632],x[2647:2640],x[2655:2648],x[2663:2656],x[2671:2664],x[2679:2672],x[2687:2680],x[2567:2560],x[2575:2568],x[2583:2576],x[2591:2584],x[2599:2592],x[2607:2600],x[2615:2608],x[2623:2616],x[2503:2496],x[2511:2504],x[2519:2512],x[2527:2520],x[2535:2528],x[2543:2536],x[2551:2544],x[2559:2552],x[2439:2432],x[2447:2440],x[2455:2448],x[2463:2456],x[2471:2464],x[2479:2472],x[2487:2480],x[2495:2488],x[2375:2368],x[2383:2376],x[2391:2384],x[2399:2392],x[2407:2400],x[2415:2408],x[2423:2416],x[2431:2424],x[2311:2304],x[2319:2312],x[2327:2320],x[2335:2328],x[2343:2336],x[2351:2344],x[2359:2352],x[2367:2360],x[2247:2240],x[2255:2248],x[2263:2256],x[2271:2264],x[2279:2272],x[2287:2280],x[2295:2288],x[2303:2296],x[2183:2176],x[2191:2184],x[2199:2192],x[2207:2200],x[2215:2208],x[2223:2216],x[2231:2224],x[2239:2232],x[2119:2112],x[2127:2120],x[2135:2128],x[2143:2136],x[2151:2144],x[2159:2152],x[2167:2160],x[2175:2168],x[2055:2048],x[2063:2056],x[2071:2064],x[2079:2072],x[2087:2080],x[2095:2088],x[2103:2096],x[2111:2104],x[1991:1984],x[1999:1992],x[2007:2000],x[2015:2008],x[2023:2016],x[2031:2024],x[2039:2032],x[2047:2040],x[1927:1920],x[1935:1928],x[1943:1936],x[1951:1944],x[1959:1952],x[1967:1960],x[1975:1968],x[1983:1976],x[1863:1856],x[1871:1864],x[1879:1872],x[1887:1880],x[1895:1888],x[1903:1896],x[1911:1904],x[1919:1912],x[1799:1792],x[1807:1800],x[1815:1808],x[1823:1816],x[1831:1824],x[1839:1832],x[1847:1840],x[1855:1848],x[1735:1728],x[1743:1736],x[1751:1744],x[1759:1752],x[1767:1760],x[1775:1768],x[1783:1776],x[1791:1784],x[1671:1664],x[1679:1672],x[1687:1680],x[1695:1688],x[1703:1696],x[1711:1704],x[1719:1712],x[1727:1720],x[1607:1600],x[1615:1608],x[1623:1616],x[1631:1624],x[1639:1632],x[1647:1640],x[1655:1648],x[1663:1656],x[1543:1536],x[1551:1544],x[1559:1552],x[1567:1560],x[1575:1568],x[1583:1576],x[1591:1584],x[1599:1592],x[1479:1472],x[1487:1480],x[1495:1488],x[1503:1496],x[1511:1504],x[1519:1512],x[1527:1520],x[1535:1528],x[1415:1408],x[1423:1416],x[1431:1424],x[1439:1432],x[1447:1440],x[1455:1448],x[1463:1456],x[1471:1464],x[1351:1344],x[1359:1352],x[1367:1360],x[1375:1368],x[1383:1376],x[1391:1384],x[1399:1392],x[1407:1400],x[1287:1280],x[1295:1288],x[1303:1296],x[1311:1304],x[1319:1312],x[1327:1320],x[1335:1328],x[1343:1336],x[1223:1216],x[1231:1224],x[1239:1232],x[1247:1240],x[1255:1248],x[1263:1256],x[1271:1264],x[1279:1272],x[1159:1152],x[1167:1160],x[1175:1168],x[1183:1176],x[1191:1184],x[1199:1192],x[1207:1200],x[1215:1208],x[1095:1088],x[1103:1096],x[1111:1104],x[1119:1112],x[1127:1120],x[1135:1128],x[1143:1136],x[1151:1144],x[1031:1024],x[1039:1032],x[1047:1040],x[1055:1048],x[1063:1056],x[1071:1064],x[1079:1072],x[1087:1080],x[967:960],x[975:968],x[983:976],x[991:984],x[999:992],x[1007:1000],x[1015:1008],x[1023:1016],x[903:896],x[911:904],x[919:912],x[927:920],x[935:928],x[943:936],x[951:944],x[959:952],x[839:832],x[847:840],x[855:848],x[863:856],x[871:864],x[879:872],x[887:880],x[895:888],x[775:768],x[783:776],x[791:784],x[799:792],x[807:800],x[815:808],x[823:816],x[831:824],x[711:704],x[719:712],x[727:720],x[735:728],x[743:736],x[751:744],x[759:752],x[767:760],x[647:640],x[655:648],x[663:656],x[671:664],x[679:672],x[687:680],x[695:688],x[703:696],x[583:576],x[591:584],x[599:592],x[607:600],x[615:608],x[623:616],x[631:624],x[639:632],x[519:512],x[527:520],x[535:528],x[543:536],x[551:544],x[559:552],x[567:560],x[575:568],x[455:448],x[463:456],x[471:464],x[479:472],x[487:480],x[495:488],x[503:496],x[511:504],x[391:384],x[399:392],x[407:400],x[415:408],x[423:416],x[431:424],x[439:432],x[447:440],x[327:320],x[335:328],x[343:336],x[351:344],x[359:352],x[367:360],x[375:368],x[383:376],x[263:256],x[271:264],x[279:272],x[287:280],x[295:288],x[303:296],x[311:304],x[319:312],x[199:192],x[207:200],x[215:208],x[223:216],x[231:224],x[239:232],x[247:240],x[255:248],x[135:128],x[143:136],x[151:144],x[159:152],x[167:160],x[175:168],x[183:176],x[191:184],x[71:64],x[79:72],x[87:80],x[95:88],x[103:96],x[111:104],x[119:112],x[127:120],x[7:0],x[15:8],x[23:16],x[31:24],x[39:32],x[47:40],x[55:48],x[63:56]}	

`define clog2_key(x)\
(x == 0) ? 0    : (x<16**1) ? 4: (x<16**2) ? 8: (x<16**3) ? 12: (x<16**4) ? 16: (x<16**5) ? 20: (x<16**6) ? 24: (x<16**7) ? 28: (x<16**8) ? 32: (x<16**9) ? 36: (x<16**10) ? 40: (x<16**11) ? 44: (x<16**12) ? 48: (x<16**13) ? 52: (x<16**14) ? 56: (x<16**15) ? 60: (x<16**16) ? 64: (x<16**17) ? 68: (x<16**18) ? 72: (x<16**19) ? 76: (x<16**20) ? 80: (x<16**21) ? 84: (x<16**22) ? 88: (x<16**23) ? 92: (x<16**24) ? 96: (x<16**25) ? 100: (x<16**26) ? 104: (x<16**27) ? 108: (x<16**28) ? 112: (x<16**29) ? 116: (x<16**30) ? 120: (x<16**31) ? 124: (x<16**32) ? 128: (x<16**33) ? 132: (x<16**34) ? 136: (x<16**35) ? 140: (x<16**36) ? 144: (x<16**37) ? 148: (x<16**38) ? 152: (x<16**39) ? 156: (x<16**40) ? 160: (x<16**41) ? 164: (x<16**42) ? 168: (x<16**43) ? 172: (x<16**44) ? 176: (x<16**45) ? 180: (x<16**46) ? 184: (x<16**47) ? 188: (x<16**48) ? 192: (x<16**49) ? 196: (x<16**50) ? 200: (x<16**51) ? 204: (x<16**52) ? 208: (x<16**53) ? 212: (x<16**54) ? 216: (x<16**55) ? 220: (x<16**56) ? 224: (x<16**57) ? 228: (x<16**58) ? 232: (x<16**59) ? 236: (x<16**60) ? 240: (x<16**61) ? 244: (x<16**62) ? 248: (x<16**63) ? 252: (x<16**64) ? 256: (x<16**65) ? 260: (x<16**66) ? 264: (x<16**67) ? 268: (x<16**68) ? 272: (x<16**69) ? 276: (x<16**70) ? 280: (x<16**71) ? 284: (x<16**72) ? 288: (x<16**73) ? 292: (x<16**74) ? 296: (x<16**75) ? 300: (x<16**76) ? 304: (x<16**77) ? 308: (x<16**78) ? 312: (x<16**79) ? 316: (x<16**80) ? 320: (x<16**81) ? 324: (x<16**82) ? 328: (x<16**83) ? 332: (x<16**84) ? 336: (x<16**85) ? 340: (x<16**86) ? 344: (x<16**87) ? 348: (x<16**88) ? 352: (x<16**89) ? 356: (x<16**90) ? 360: (x<16**91) ? 364: (x<16**92) ? 368: (x<16**93) ? 372: (x<16**94) ? 376: (x<16**95) ? 380: (x<16**96) ? 384: (x<16**97) ? 388: (x<16**98) ? 392: (x<16**99) ? 396: (x<16**100) ? 400: (x<16**101) ? 404: (x<16**102) ? 408: (x<16**103) ? 412: (x<16**104) ? 416: (x<16**105) ? 420: (x<16**106) ? 424: (x<16**107) ? 428: (x<16**108) ? 432: (x<16**109) ? 436: (x<16**110) ? 440: (x<16**111) ? 444: (x<16**112) ? 448: (x<16**113) ? 452: (x<16**114) ? 456: (x<16**115) ? 460: (x<16**116) ? 464: (x<16**117) ? 468: (x<16**118) ? 472: (x<16**119) ? 476: (x<16**120) ? 480: (x<16**121) ? 484: (x<16**122) ? 488: (x<16**123) ? 492: (x<16**124) ? 496: (x<16**125) ? 500: (x<16**126) ? 504: (x<16**127) ? 508: (x<16**128) ? 512 : -1

`define rotate_key(x)\
{x[455:448],x[463:456],x[471:464],x[479:472],x[487:480],x[495:488],x[503:496],x[511:504],x[391:384],x[399:392],x[407:400],x[415:408],x[423:416],x[431:424],x[439:432],x[447:440],x[327:320],x[335:328],x[343:336],x[351:344],x[359:352],x[367:360],x[375:368],x[383:376],x[263:256],x[271:264],x[279:272],x[287:280],x[295:288],x[303:296],x[311:304],x[319:312],x[199:192],x[207:200],x[215:208],x[223:216],x[231:224],x[239:232],x[247:240],x[255:248],x[135:128],x[143:136],x[151:144],x[159:152],x[167:160],x[175:168],x[183:176],x[191:184],x[71:64],x[79:72],x[87:80],x[95:88],x[103:96],x[111:104],x[119:112],x[127:120],x[7:0],x[15:8],x[23:16],x[31:24],x[39:32],x[47:40],x[55:48],x[63:56]}	

`define rotate_D(x)\
{x[63:0],x[127:64],x[191:128],x[255:192]}

// Massage example 2 
`define M1		64'h1122334455667711
`define M2		64'h2233445566771122
`define M3		64'h3344556677112233
`define M4		64'h4455667711223344
`define M5		64'h5566771122334455
`define M6		64'h6677112233445566
`define M7		64'h7711223344556677

`define M_array_2  {`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1}

// Massage example 3 

`define M_array_3  {`M2,	 `M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1,	`M7,	`M6,	`M5,	`M4,	`M3,	`M2,	`M1}
