`include "parameters.vh"
//
//This module is responsible for the computation of 16 steps (16 words) itself.
//We have designed it in such a way that we would not have to use a clock in order to save FF resources
//
//
module A_computation_loop      
( 
    input  wire 		         		clk,
	input  wire 		          		reset,
	input  wire 				   		enable,
	input  wire  [11:0] 		  		r,
    input  wire  [168*`w-1:0]   		S, 
	input  wire  [16*`b-1:0]			R_shift,
	input  wire  [16*`b-1:0]    		L_shift,
	input  wire  [`n*`w-1:0] 			A,
	output reg   						N_to_A_en,
	output reg 							iterative_en,
	output wire  [11:0]			  		A_round_i,
    output wire  [`c*`w-1:0]    		A_steps,
	output reg 				  			done,
	output reg 							A_shift_stop
             
	
);

	reg [11:0]					j = 0	 ; // rounds index 
	reg [2:0]			    	state = 0;                 

always @ (posedge clk) 	
begin
	if (reset)
	begin
		state <= 0;
		j <= 0;	
		done <= 0;
		A_shift_stop <= 1;
		N_to_A_en <= 0;
		iterative_en <=0;
	end
	else
	begin
		case (state)
			0:
			begin
			if (enable)
				state <= 1;
				done <= 0;
				j <= 0;
			end
			1:
			begin
			N_to_A_en <= 1;
			A_shift_stop <= 0;
			state <= 2;
			end
			2:
			begin
			iterative_en <=1;
			state <=3;
			end
			3:
			begin
				N_to_A_en <= 0;
				iterative_en <=0;
				if ((j < r) && enable)
				begin		
					j <= j + 1;	
				end
				else 			// end of cf indecator
				begin
					done <= 1;
					state <= 4;
				end
				if(j==(r-1))
					A_shift_stop <= 1;		
			end	
			4:
			begin
			end
		endcase
	end
end


assign A_round_i = j; 


// MD6 16 steps, every round 
	assign A_steps[0 *`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(0 )*`w+:`w]   ^ A[((`n + 0) -  `t0 )*`w+:`w])^((A[(`n + 0 -  `t1 )*`w+:`w]  & A[(`n + 0 -  `t2 )*`w+:`w])  ^ (A[(`n + 0 -  `t3 )*`w+:`w]  & A[(`n + 0 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(0 )*`w+:`w]   ^ A[((`n + 0) -  `t0 )*`w+:`w])^((A[(`n + 0 -  `t1 )*`w+:`w]  & A[(`n + 0 -  `t2 )*`w+:`w])  ^ (A[(`n + 0 -  `t3 )*`w+:`w]  & A[(`n + 0 -  `t4 )*`w+:`w])))) >> R_shift[1 *`b-1: 0* `b])))^((((((S[(j)*`w+:`w] ^ A[(0 )*`w+:`w]   ^ A[((`n + 0) -  `t0 )*`w+:`w])^((A[(`n + 0 -  `t1 )*`w+:`w]  & A[(`n + 0 -  `t2 )*`w+:`w])  ^ (A[(`n + 0 -  `t3 )*`w+:`w]  & A[(`n + 0 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(0 )*`w+:`w]   ^ A[((`n + 0) -  `t0 )*`w+:`w])^((A[(`n + 0 -  `t1 )*`w+:`w]  & A[(`n + 0 -  `t2 )*`w+:`w])  ^ (A[(`n + 0 -  `t3 )*`w+:`w]  & A[(`n + 0 -  `t4 )*`w+:`w])))) >> R_shift[1 *`b-1: 0* `b])))) << L_shift[1 *`b-1:0 *`b]));
	assign A_steps[1 *`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(1 )*`w+:`w]   ^ A[((`n + 1) -  `t0 )*`w+:`w])^((A[(`n + 1 -  `t1 )*`w+:`w]  & A[(`n + 1 -  `t2 )*`w+:`w])  ^ (A[(`n + 1 -  `t3 )*`w+:`w]  & A[(`n + 1 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(1 )*`w+:`w]   ^ A[((`n + 1) -  `t0 )*`w+:`w])^((A[(`n + 1 -  `t1 )*`w+:`w]  & A[(`n + 1 -  `t2 )*`w+:`w])  ^ (A[(`n + 1 -  `t3 )*`w+:`w]  & A[(`n + 1 -  `t4 )*`w+:`w])))) >> R_shift[2 *`b-1: 1* `b])))^((((((S[(j)*`w+:`w] ^ A[(1 )*`w+:`w]   ^ A[((`n + 1) -  `t0 )*`w+:`w])^((A[(`n + 1 -  `t1 )*`w+:`w]  & A[(`n + 1 -  `t2 )*`w+:`w])  ^ (A[(`n + 1 -  `t3 )*`w+:`w]  & A[(`n + 1 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(1 )*`w+:`w]   ^ A[((`n + 1) -  `t0 )*`w+:`w])^((A[(`n + 1 -  `t1 )*`w+:`w]  & A[(`n + 1 -  `t2 )*`w+:`w])  ^ (A[(`n + 1 -  `t3 )*`w+:`w]  & A[(`n + 1 -  `t4 )*`w+:`w])))) >> R_shift[2 *`b-1: 1* `b])))) << L_shift[2 *`b-1:1 *`b]));
	assign A_steps[2 *`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(2 )*`w+:`w]   ^ A[((`n + 2) -  `t0 )*`w+:`w])^((A[(`n + 2 -  `t1 )*`w+:`w]  & A[(`n + 2 -  `t2 )*`w+:`w])  ^ (A[(`n + 2 -  `t3 )*`w+:`w]  & A[(`n + 2 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(2 )*`w+:`w]   ^ A[((`n + 2) -  `t0 )*`w+:`w])^((A[(`n + 2 -  `t1 )*`w+:`w]  & A[(`n + 2 -  `t2 )*`w+:`w])  ^ (A[(`n + 2 -  `t3 )*`w+:`w]  & A[(`n + 2 -  `t4 )*`w+:`w])))) >> R_shift[3 *`b-1: 2* `b])))^((((((S[(j)*`w+:`w] ^ A[(2 )*`w+:`w]   ^ A[((`n + 2) -  `t0 )*`w+:`w])^((A[(`n + 2 -  `t1 )*`w+:`w]  & A[(`n + 2 -  `t2 )*`w+:`w])  ^ (A[(`n + 2 -  `t3 )*`w+:`w]  & A[(`n + 2 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(2 )*`w+:`w]   ^ A[((`n + 2) -  `t0 )*`w+:`w])^((A[(`n + 2 -  `t1 )*`w+:`w]  & A[(`n + 2 -  `t2 )*`w+:`w])  ^ (A[(`n + 2 -  `t3 )*`w+:`w]  & A[(`n + 2 -  `t4 )*`w+:`w])))) >> R_shift[3 *`b-1: 2* `b])))) << L_shift[3 *`b-1:2 *`b]));
	assign A_steps[3 *`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(3 )*`w+:`w]   ^ A[((`n + 3) -  `t0 )*`w+:`w])^((A[(`n + 3 -  `t1 )*`w+:`w]  & A[(`n + 3 -  `t2 )*`w+:`w])  ^ (A[(`n + 3 -  `t3 )*`w+:`w]  & A[(`n + 3 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(3 )*`w+:`w]   ^ A[((`n + 3) -  `t0 )*`w+:`w])^((A[(`n + 3 -  `t1 )*`w+:`w]  & A[(`n + 3 -  `t2 )*`w+:`w])  ^ (A[(`n + 3 -  `t3 )*`w+:`w]  & A[(`n + 3 -  `t4 )*`w+:`w])))) >> R_shift[4 *`b-1: 3* `b])))^((((((S[(j)*`w+:`w] ^ A[(3 )*`w+:`w]   ^ A[((`n + 3) -  `t0 )*`w+:`w])^((A[(`n + 3 -  `t1 )*`w+:`w]  & A[(`n + 3 -  `t2 )*`w+:`w])  ^ (A[(`n + 3 -  `t3 )*`w+:`w]  & A[(`n + 3 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(3 )*`w+:`w]   ^ A[((`n + 3) -  `t0 )*`w+:`w])^((A[(`n + 3 -  `t1 )*`w+:`w]  & A[(`n + 3 -  `t2 )*`w+:`w])  ^ (A[(`n + 3 -  `t3 )*`w+:`w]  & A[(`n + 3 -  `t4 )*`w+:`w])))) >> R_shift[4 *`b-1: 3* `b])))) << L_shift[4 *`b-1:3 *`b]));
	assign A_steps[4 *`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(4 )*`w+:`w]   ^ A[((`n + 4) -  `t0 )*`w+:`w])^((A[(`n + 4 -  `t1 )*`w+:`w]  & A[(`n + 4 -  `t2 )*`w+:`w])  ^ (A[(`n + 4 -  `t3 )*`w+:`w]  & A[(`n + 4 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(4 )*`w+:`w]   ^ A[((`n + 4) -  `t0 )*`w+:`w])^((A[(`n + 4 -  `t1 )*`w+:`w]  & A[(`n + 4 -  `t2 )*`w+:`w])  ^ (A[(`n + 4 -  `t3 )*`w+:`w]  & A[(`n + 4 -  `t4 )*`w+:`w])))) >> R_shift[5 *`b-1: 4* `b])))^((((((S[(j)*`w+:`w] ^ A[(4 )*`w+:`w]   ^ A[((`n + 4) -  `t0 )*`w+:`w])^((A[(`n + 4 -  `t1 )*`w+:`w]  & A[(`n + 4 -  `t2 )*`w+:`w])  ^ (A[(`n + 4 -  `t3 )*`w+:`w]  & A[(`n + 4 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(4 )*`w+:`w]   ^ A[((`n + 4) -  `t0 )*`w+:`w])^((A[(`n + 4 -  `t1 )*`w+:`w]  & A[(`n + 4 -  `t2 )*`w+:`w])  ^ (A[(`n + 4 -  `t3 )*`w+:`w]  & A[(`n + 4 -  `t4 )*`w+:`w])))) >> R_shift[5 *`b-1: 4* `b])))) << L_shift[5 *`b-1:4 *`b]));
	assign A_steps[5 *`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(5 )*`w+:`w]   ^ A[((`n + 5) -  `t0 )*`w+:`w])^((A[(`n + 5 -  `t1 )*`w+:`w]  & A[(`n + 5 -  `t2 )*`w+:`w])  ^ (A[(`n + 5 -  `t3 )*`w+:`w]  & A[(`n + 5 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(5 )*`w+:`w]   ^ A[((`n + 5) -  `t0 )*`w+:`w])^((A[(`n + 5 -  `t1 )*`w+:`w]  & A[(`n + 5 -  `t2 )*`w+:`w])  ^ (A[(`n + 5 -  `t3 )*`w+:`w]  & A[(`n + 5 -  `t4 )*`w+:`w])))) >> R_shift[6 *`b-1: 5* `b])))^((((((S[(j)*`w+:`w] ^ A[(5 )*`w+:`w]   ^ A[((`n + 5) -  `t0 )*`w+:`w])^((A[(`n + 5 -  `t1 )*`w+:`w]  & A[(`n + 5 -  `t2 )*`w+:`w])  ^ (A[(`n + 5 -  `t3 )*`w+:`w]  & A[(`n + 5 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(5 )*`w+:`w]   ^ A[((`n + 5) -  `t0 )*`w+:`w])^((A[(`n + 5 -  `t1 )*`w+:`w]  & A[(`n + 5 -  `t2 )*`w+:`w])  ^ (A[(`n + 5 -  `t3 )*`w+:`w]  & A[(`n + 5 -  `t4 )*`w+:`w])))) >> R_shift[6 *`b-1: 5* `b])))) << L_shift[6 *`b-1:5 *`b]));
	assign A_steps[6 *`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(6 )*`w+:`w]   ^ A[((`n + 6) -  `t0 )*`w+:`w])^((A[(`n + 6 -  `t1 )*`w+:`w]  & A[(`n + 6 -  `t2 )*`w+:`w])  ^ (A[(`n + 6 -  `t3 )*`w+:`w]  & A[(`n + 6 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(6 )*`w+:`w]   ^ A[((`n + 6) -  `t0 )*`w+:`w])^((A[(`n + 6 -  `t1 )*`w+:`w]  & A[(`n + 6 -  `t2 )*`w+:`w])  ^ (A[(`n + 6 -  `t3 )*`w+:`w]  & A[(`n + 6 -  `t4 )*`w+:`w])))) >> R_shift[7 *`b-1: 6* `b])))^((((((S[(j)*`w+:`w] ^ A[(6 )*`w+:`w]   ^ A[((`n + 6) -  `t0 )*`w+:`w])^((A[(`n + 6 -  `t1 )*`w+:`w]  & A[(`n + 6 -  `t2 )*`w+:`w])  ^ (A[(`n + 6 -  `t3 )*`w+:`w]  & A[(`n + 6 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(6 )*`w+:`w]   ^ A[((`n + 6) -  `t0 )*`w+:`w])^((A[(`n + 6 -  `t1 )*`w+:`w]  & A[(`n + 6 -  `t2 )*`w+:`w])  ^ (A[(`n + 6 -  `t3 )*`w+:`w]  & A[(`n + 6 -  `t4 )*`w+:`w])))) >> R_shift[7 *`b-1: 6* `b])))) << L_shift[7 *`b-1:6 *`b]));
	assign A_steps[7 *`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(7 )*`w+:`w]   ^ A[((`n + 7) -  `t0 )*`w+:`w])^((A[(`n + 7 -  `t1 )*`w+:`w]  & A[(`n + 7 -  `t2 )*`w+:`w])  ^ (A[(`n + 7 -  `t3 )*`w+:`w]  & A[(`n + 7 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(7 )*`w+:`w]   ^ A[((`n + 7) -  `t0 )*`w+:`w])^((A[(`n + 7 -  `t1 )*`w+:`w]  & A[(`n + 7 -  `t2 )*`w+:`w])  ^ (A[(`n + 7 -  `t3 )*`w+:`w]  & A[(`n + 7 -  `t4 )*`w+:`w])))) >> R_shift[8 *`b-1: 7* `b])))^((((((S[(j)*`w+:`w] ^ A[(7 )*`w+:`w]   ^ A[((`n + 7) -  `t0 )*`w+:`w])^((A[(`n + 7 -  `t1 )*`w+:`w]  & A[(`n + 7 -  `t2 )*`w+:`w])  ^ (A[(`n + 7 -  `t3 )*`w+:`w]  & A[(`n + 7 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(7 )*`w+:`w]   ^ A[((`n + 7) -  `t0 )*`w+:`w])^((A[(`n + 7 -  `t1 )*`w+:`w]  & A[(`n + 7 -  `t2 )*`w+:`w])  ^ (A[(`n + 7 -  `t3 )*`w+:`w]  & A[(`n + 7 -  `t4 )*`w+:`w])))) >> R_shift[8 *`b-1: 7* `b])))) << L_shift[8 *`b-1:7 *`b]));
	assign A_steps[8 *`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(8 )*`w+:`w]   ^ A[((`n + 8) -  `t0 )*`w+:`w])^((A[(`n + 8 -  `t1 )*`w+:`w]  & A[(`n + 8 -  `t2 )*`w+:`w])  ^ (A[(`n + 8 -  `t3 )*`w+:`w]  & A[(`n + 8 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(8 )*`w+:`w]   ^ A[((`n + 8) -  `t0 )*`w+:`w])^((A[(`n + 8 -  `t1 )*`w+:`w]  & A[(`n + 8 -  `t2 )*`w+:`w])  ^ (A[(`n + 8 -  `t3 )*`w+:`w]  & A[(`n + 8 -  `t4 )*`w+:`w])))) >> R_shift[9 *`b-1: 8* `b])))^((((((S[(j)*`w+:`w] ^ A[(8 )*`w+:`w]   ^ A[((`n + 8) -  `t0 )*`w+:`w])^((A[(`n + 8 -  `t1 )*`w+:`w]  & A[(`n + 8 -  `t2 )*`w+:`w])  ^ (A[(`n + 8 -  `t3 )*`w+:`w]  & A[(`n + 8 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(8 )*`w+:`w]   ^ A[((`n + 8) -  `t0 )*`w+:`w])^((A[(`n + 8 -  `t1 )*`w+:`w]  & A[(`n + 8 -  `t2 )*`w+:`w])  ^ (A[(`n + 8 -  `t3 )*`w+:`w]  & A[(`n + 8 -  `t4 )*`w+:`w])))) >> R_shift[9 *`b-1: 8* `b])))) << L_shift[9 *`b-1:8 *`b]));
	assign A_steps[9 *`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(9 )*`w+:`w]   ^ A[((`n + 9) -  `t0 )*`w+:`w])^((A[(`n + 9 -  `t1 )*`w+:`w]  & A[(`n + 9 -  `t2 )*`w+:`w])  ^ (A[(`n + 9 -  `t3 )*`w+:`w]  & A[(`n + 9 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(9 )*`w+:`w]   ^ A[((`n + 9) -  `t0 )*`w+:`w])^((A[(`n + 9 -  `t1 )*`w+:`w]  & A[(`n + 9 -  `t2 )*`w+:`w])  ^ (A[(`n + 9 -  `t3 )*`w+:`w]  & A[(`n + 9 -  `t4 )*`w+:`w])))) >> R_shift[10*`b-1: 9* `b])))^((((((S[(j)*`w+:`w] ^ A[(9 )*`w+:`w]   ^ A[((`n + 9) -  `t0 )*`w+:`w])^((A[(`n + 9 -  `t1 )*`w+:`w]  & A[(`n + 9 -  `t2 )*`w+:`w])  ^ (A[(`n + 9 -  `t3 )*`w+:`w]  & A[(`n + 9 -  `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(9 )*`w+:`w]   ^ A[((`n + 9) -  `t0 )*`w+:`w])^((A[(`n + 9 -  `t1 )*`w+:`w]  & A[(`n + 9 -  `t2 )*`w+:`w])  ^ (A[(`n + 9 -  `t3 )*`w+:`w]  & A[(`n + 9 -  `t4 )*`w+:`w])))) >> R_shift[10*`b-1: 9* `b])))) << L_shift[10*`b-1:9 *`b]));
	assign A_steps[10*`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(10 )*`w+:`w]  ^ A[((`n + 10) - `t0 )*`w+:`w])^((A[(`n + 10 - `t1 )*`w+:`w]  & A[(`n + 10 - `t2 )*`w+:`w])  ^ (A[(`n + 10 - `t3 )*`w+:`w]  & A[(`n + 10 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(10 )*`w+:`w]  ^ A[((`n + 10) - `t0 )*`w+:`w])^((A[(`n + 10 - `t1 )*`w+:`w]  & A[(`n + 10 - `t2 )*`w+:`w])  ^ (A[(`n + 10 - `t3 )*`w+:`w]  & A[(`n + 10 - `t4 )*`w+:`w])))) >> R_shift[11*`b-1: 10*`b])))^((((((S[(j)*`w+:`w] ^ A[(10 )*`w+:`w]  ^ A[((`n + 10) - `t0 )*`w+:`w])^((A[(`n + 10 - `t1 )*`w+:`w]  & A[(`n + 10 - `t2 )*`w+:`w])  ^ (A[(`n + 10 - `t3 )*`w+:`w]  & A[(`n + 10 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(10 )*`w+:`w]  ^ A[((`n + 10) - `t0 )*`w+:`w])^((A[(`n + 10 - `t1 )*`w+:`w]  & A[(`n + 10 - `t2 )*`w+:`w])  ^ (A[(`n + 10 - `t3 )*`w+:`w]  & A[(`n + 10 - `t4 )*`w+:`w])))) >> R_shift[11*`b-1: 10*`b])))) << L_shift[11*`b-1:10*`b]));
	assign A_steps[11*`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(11 )*`w+:`w]  ^ A[((`n + 11) - `t0 )*`w+:`w])^((A[(`n + 11 - `t1 )*`w+:`w]  & A[(`n + 11 - `t2 )*`w+:`w])  ^ (A[(`n + 11 - `t3 )*`w+:`w]  & A[(`n + 11 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(11 )*`w+:`w]  ^ A[((`n + 11) - `t0 )*`w+:`w])^((A[(`n + 11 - `t1 )*`w+:`w]  & A[(`n + 11 - `t2 )*`w+:`w])  ^ (A[(`n + 11 - `t3 )*`w+:`w]  & A[(`n + 11 - `t4 )*`w+:`w])))) >> R_shift[12*`b-1: 11*`b])))^((((((S[(j)*`w+:`w] ^ A[(11 )*`w+:`w]  ^ A[((`n + 11) - `t0 )*`w+:`w])^((A[(`n + 11 - `t1 )*`w+:`w]  & A[(`n + 11 - `t2 )*`w+:`w])  ^ (A[(`n + 11 - `t3 )*`w+:`w]  & A[(`n + 11 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(11 )*`w+:`w]  ^ A[((`n + 11) - `t0 )*`w+:`w])^((A[(`n + 11 - `t1 )*`w+:`w]  & A[(`n + 11 - `t2 )*`w+:`w])  ^ (A[(`n + 11 - `t3 )*`w+:`w]  & A[(`n + 11 - `t4 )*`w+:`w])))) >> R_shift[12*`b-1: 11*`b])))) << L_shift[12*`b-1:11*`b]));
	assign A_steps[12*`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(12 )*`w+:`w]  ^ A[((`n + 12) - `t0 )*`w+:`w])^((A[(`n + 12 - `t1 )*`w+:`w]  & A[(`n + 12 - `t2 )*`w+:`w])  ^ (A[(`n + 12 - `t3 )*`w+:`w]  & A[(`n + 12 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(12 )*`w+:`w]  ^ A[((`n + 12) - `t0 )*`w+:`w])^((A[(`n + 12 - `t1 )*`w+:`w]  & A[(`n + 12 - `t2 )*`w+:`w])  ^ (A[(`n + 12 - `t3 )*`w+:`w]  & A[(`n + 12 - `t4 )*`w+:`w])))) >> R_shift[13*`b-1: 12*`b])))^((((((S[(j)*`w+:`w] ^ A[(12 )*`w+:`w]  ^ A[((`n + 12) - `t0 )*`w+:`w])^((A[(`n + 12 - `t1 )*`w+:`w]  & A[(`n + 12 - `t2 )*`w+:`w])  ^ (A[(`n + 12 - `t3 )*`w+:`w]  & A[(`n + 12 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(12 )*`w+:`w]  ^ A[((`n + 12) - `t0 )*`w+:`w])^((A[(`n + 12 - `t1 )*`w+:`w]  & A[(`n + 12 - `t2 )*`w+:`w])  ^ (A[(`n + 12 - `t3 )*`w+:`w]  & A[(`n + 12 - `t4 )*`w+:`w])))) >> R_shift[13*`b-1: 12*`b])))) << L_shift[13*`b-1:12*`b]));
	assign A_steps[13*`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(13 )*`w+:`w]  ^ A[((`n + 13) - `t0 )*`w+:`w])^((A[(`n + 13 - `t1 )*`w+:`w]  & A[(`n + 13 - `t2 )*`w+:`w])  ^ (A[(`n + 13 - `t3 )*`w+:`w]  & A[(`n + 13 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(13 )*`w+:`w]  ^ A[((`n + 13) - `t0 )*`w+:`w])^((A[(`n + 13 - `t1 )*`w+:`w]  & A[(`n + 13 - `t2 )*`w+:`w])  ^ (A[(`n + 13 - `t3 )*`w+:`w]  & A[(`n + 13 - `t4 )*`w+:`w])))) >> R_shift[14*`b-1: 13*`b])))^((((((S[(j)*`w+:`w] ^ A[(13 )*`w+:`w]  ^ A[((`n + 13) - `t0 )*`w+:`w])^((A[(`n + 13 - `t1 )*`w+:`w]  & A[(`n + 13 - `t2 )*`w+:`w])  ^ (A[(`n + 13 - `t3 )*`w+:`w]  & A[(`n + 13 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(13 )*`w+:`w]  ^ A[((`n + 13) - `t0 )*`w+:`w])^((A[(`n + 13 - `t1 )*`w+:`w]  & A[(`n + 13 - `t2 )*`w+:`w])  ^ (A[(`n + 13 - `t3 )*`w+:`w]  & A[(`n + 13 - `t4 )*`w+:`w])))) >> R_shift[14*`b-1: 13*`b])))) << L_shift[14*`b-1:13*`b]));
	assign A_steps[14*`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(14 )*`w+:`w]  ^ A[((`n + 14) - `t0 )*`w+:`w])^((A[(`n + 14 - `t1 )*`w+:`w]  & A[(`n + 14 - `t2 )*`w+:`w])  ^ (A[(`n + 14 - `t3 )*`w+:`w]  & A[(`n + 14 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(14 )*`w+:`w]  ^ A[((`n + 14) - `t0 )*`w+:`w])^((A[(`n + 14 - `t1 )*`w+:`w]  & A[(`n + 14 - `t2 )*`w+:`w])  ^ (A[(`n + 14 - `t3 )*`w+:`w]  & A[(`n + 14 - `t4 )*`w+:`w])))) >> R_shift[15*`b-1: 14*`b])))^((((((S[(j)*`w+:`w] ^ A[(14 )*`w+:`w]  ^ A[((`n + 14) - `t0 )*`w+:`w])^((A[(`n + 14 - `t1 )*`w+:`w]  & A[(`n + 14 - `t2 )*`w+:`w])  ^ (A[(`n + 14 - `t3 )*`w+:`w]  & A[(`n + 14 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(14 )*`w+:`w]  ^ A[((`n + 14) - `t0 )*`w+:`w])^((A[(`n + 14 - `t1 )*`w+:`w]  & A[(`n + 14 - `t2 )*`w+:`w])  ^ (A[(`n + 14 - `t3 )*`w+:`w]  & A[(`n + 14 - `t4 )*`w+:`w])))) >> R_shift[15*`b-1: 14*`b])))) << L_shift[15*`b-1:14*`b]));
	assign A_steps[15*`w+:`w]  =  (((S[(j)*`w+:`w] ^ A[(15 )*`w+:`w]  ^ A[((`n + 15) - `t0 )*`w+:`w])^((A[(`n + 15 - `t1 )*`w+:`w]  & A[(`n + 15 - `t2 )*`w+:`w])  ^ (A[(`n + 15 - `t3 )*`w+:`w]  & A[(`n + 15 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(15 )*`w+:`w]  ^ A[((`n + 15) - `t0 )*`w+:`w])^((A[(`n + 15 - `t1 )*`w+:`w]  & A[(`n + 15 - `t2 )*`w+:`w])  ^ (A[(`n + 15 - `t3 )*`w+:`w]  & A[(`n + 15 - `t4 )*`w+:`w])))) >> R_shift[16*`b-1: 15*`b])))^((((((S[(j)*`w+:`w] ^ A[(15 )*`w+:`w]  ^ A[((`n + 15) - `t0 )*`w+:`w])^((A[(`n + 15 - `t1 )*`w+:`w]  & A[(`n + 15 - `t2 )*`w+:`w])  ^ (A[(`n + 15 - `t3 )*`w+:`w]  & A[(`n + 15 - `t4 )*`w+:`w])))^(((((S[(j)*`w+:`w] ^ A[(15 )*`w+:`w]  ^ A[((`n + 15) - `t0 )*`w+:`w])^((A[(`n + 15 - `t1 )*`w+:`w]  & A[(`n + 15 - `t2 )*`w+:`w])  ^ (A[(`n + 15 - `t3 )*`w+:`w]  & A[(`n + 15 - `t4 )*`w+:`w])))) >> R_shift[16*`b-1: 15*`b])))) << L_shift[16*`b-1:15*`b]));


endmodule